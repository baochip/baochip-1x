// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

`resetall
`timescale 1ns / 1ps
`default_nettype none

module memory_AesZknPlugin_rom_storage_Rom_1rs #(
    parameter wordCount = 512,
    parameter wordWidth = 32,
    parameter technology = "auto", // not used
    parameter addrWidth = $clog2(wordCount)
)
(
    input  wire                             clk,
    input  wire                             en,
    input  wire [addrWidth - 1:0]           addr,
    output reg  [wordWidth - 1:0]           data,
    input  wire                             CMBIST, // dummy pins for test insertion
    input  wire                             CMATPG, // dummy pins for test insertion
    input  wire [2:0]                       sramtrm // dummy pins for SRAM trim
);

always @(posedge clk) begin
    if (en) begin
        case (addr)
            'd0: data <= 32'b01010010101001011100011001100011;
            'd1: data <= 32'b00001001100001001111100001111100;
            'd2: data <= 32'b01101010100110011110111001110111;
            'd3: data <= 32'b11010101100011011111011001111011;
            'd4: data <= 32'b00110000000011011111111111110010;
            'd5: data <= 32'b00110110101111011101011001101011;
            'd6: data <= 32'b10100101101100011101111001101111;
            'd7: data <= 32'b00111000010101001001000111000101;
            'd8: data <= 32'b10111111010100000110000000110000;
            'd9: data <= 32'b01000000000000110000001000000001;
            'd10: data <= 32'b10100011101010011100111001100111;
            'd11: data <= 32'b10011110011111010101011000101011;
            'd12: data <= 32'b10000001000110011110011111111110;
            'd13: data <= 32'b11110011011000101011010111010111;
            'd14: data <= 32'b11010111111001100100110110101011;
            'd15: data <= 32'b11111011100110101110110001110110;
            'd16: data <= 32'b01111100010001011000111111001010;
            'd17: data <= 32'b11100011100111010001111110000010;
            'd18: data <= 32'b00111001010000001000100111001001;
            'd19: data <= 32'b10000010100001111111101001111101;
            'd20: data <= 32'b10011011000101011110111111111010;
            'd21: data <= 32'b00101111111010111011001001011001;
            'd22: data <= 32'b11111111110010011000111001000111;
            'd23: data <= 32'b10000111000010111111101111110000;
            'd24: data <= 32'b00110100111011000100000110101101;
            'd25: data <= 32'b10001110011001111011001111010100;
            'd26: data <= 32'b01000011111111010101111110100010;
            'd27: data <= 32'b01000100111010100100010110101111;
            'd28: data <= 32'b11000100101111110010001110011100;
            'd29: data <= 32'b11011110111101110101001110100100;
            'd30: data <= 32'b11101001100101101110010001110010;
            'd31: data <= 32'b11001011010110111001101111000000;
            'd32: data <= 32'b01010100110000100111010110110111;
            'd33: data <= 32'b01111011000111001110000111111101;
            'd34: data <= 32'b10010100101011100011110110010011;
            'd35: data <= 32'b00110010011010100100110000100110;
            'd36: data <= 32'b10100110010110100110110000110110;
            'd37: data <= 32'b11000010010000010111111000111111;
            'd38: data <= 32'b00100011000000101111010111110111;
            'd39: data <= 32'b00111101010011111000001111001100;
            'd40: data <= 32'b11101110010111000110100000110100;
            'd41: data <= 32'b01001100111101000101000110100101;
            'd42: data <= 32'b10010101001101001101000111100101;
            'd43: data <= 32'b00001011000010001111100111110001;
            'd44: data <= 32'b01000010100100111110001001110001;
            'd45: data <= 32'b11111010011100111010101111011000;
            'd46: data <= 32'b11000011010100110110001000110001;
            'd47: data <= 32'b01001110001111110010101000010101;
            'd48: data <= 32'b00001000000011000000100000000100;
            'd49: data <= 32'b00101110010100101001010111000111;
            'd50: data <= 32'b10100001011001010100011000100011;
            'd51: data <= 32'b01100110010111101001110111000011;
            'd52: data <= 32'b00101000001010000011000000011000;
            'd53: data <= 32'b11011001101000010011011110010110;
            'd54: data <= 32'b00100100000011110000101000000101;
            'd55: data <= 32'b10110010101101010010111110011010;
            'd56: data <= 32'b01110110000010010000111000000111;
            'd57: data <= 32'b01011011001101100010010000010010;
            'd58: data <= 32'b10100010100110110001101110000000;
            'd59: data <= 32'b01001001001111011101111111100010;
            'd60: data <= 32'b01101101001001101100110111101011;
            'd61: data <= 32'b10001011011010010100111000100111;
            'd62: data <= 32'b11010001110011010111111110110010;
            'd63: data <= 32'b00100101100111111110101001110101;
            'd64: data <= 32'b01110010000110110001001000001001;
            'd65: data <= 32'b11111000100111100001110110000011;
            'd66: data <= 32'b11110110011101000101100000101100;
            'd67: data <= 32'b01100100001011100011010000011010;
            'd68: data <= 32'b10000110001011010011011000011011;
            'd69: data <= 32'b01101000101100101101110001101110;
            'd70: data <= 32'b10011000111011101011010001011010;
            'd71: data <= 32'b00010110111110110101101110100000;
            'd72: data <= 32'b11010100111101101010010001010010;
            'd73: data <= 32'b10100100010011010111011000111011;
            'd74: data <= 32'b01011100011000011011011111010110;
            'd75: data <= 32'b11001100110011100111110110110011;
            'd76: data <= 32'b01011101011110110101001000101001;
            'd77: data <= 32'b01100101001111101101110111100011;
            'd78: data <= 32'b10110110011100010101111000101111;
            'd79: data <= 32'b10010010100101110001001110000100;
            'd80: data <= 32'b01101100111101011010011001010011;
            'd81: data <= 32'b01110000011010001011100111010001;
            'd82: data <= 32'b01001000000000000000000000000000;
            'd83: data <= 32'b01010000001011001100000111101101;
            'd84: data <= 32'b11111101011000000100000000100000;
            'd85: data <= 32'b11101101000111111110001111111100;
            'd86: data <= 32'b10111001110010000111100110110001;
            'd87: data <= 32'b11011010111011011011011001011011;
            'd88: data <= 32'b01011110101111101101010001101010;
            'd89: data <= 32'b00010101010001101000110111001011;
            'd90: data <= 32'b01000110110110010110011110111110;
            'd91: data <= 32'b01010111010010110111001000111001;
            'd92: data <= 32'b10100111110111101001010001001010;
            'd93: data <= 32'b10001101110101001001100001001100;
            'd94: data <= 32'b10011101111010001011000001011000;
            'd95: data <= 32'b10000100010010101000010111001111;
            'd96: data <= 32'b10010000011010111011101111010000;
            'd97: data <= 32'b11011000001010101100010111101111;
            'd98: data <= 32'b10101011111001010100111110101010;
            'd99: data <= 32'b00000000000101101110110111111011;
            'd100: data <= 32'b10001100110001011000011001000011;
            'd101: data <= 32'b10111100110101111001101001001101;
            'd102: data <= 32'b11010011010101010110011000110011;
            'd103: data <= 32'b00001010100101000001000110000101;
            'd104: data <= 32'b11110111110011111000101001000101;
            'd105: data <= 32'b11100100000100001110100111111001;
            'd106: data <= 32'b01011000000001100000010000000010;
            'd107: data <= 32'b00000101100000011111111001111111;
            'd108: data <= 32'b10111000111100001010000001010000;
            'd109: data <= 32'b10110011010001000111100000111100;
            'd110: data <= 32'b01000101101110100010010110011111;
            'd111: data <= 32'b00000110111000110100101110101000;
            'd112: data <= 32'b11010000111100111010001001010001;
            'd113: data <= 32'b00101100111111100101110110100011;
            'd114: data <= 32'b00011110110000001000000001000000;
            'd115: data <= 32'b10001111100010100000010110001111;
            'd116: data <= 32'b11001010101011010011111110010010;
            'd117: data <= 32'b00111111101111000010000110011101;
            'd118: data <= 32'b00001111010010000111000000111000;
            'd119: data <= 32'b00000010000001001111000111110101;
            'd120: data <= 32'b11000001110111110110001110111100;
            'd121: data <= 32'b10101111110000010111011110110110;
            'd122: data <= 32'b10111101011101011010111111011010;
            'd123: data <= 32'b00000011011000110100001000100001;
            'd124: data <= 32'b00000001001100000010000000010000;
            'd125: data <= 32'b00010011000110101110010111111111;
            'd126: data <= 32'b10001010000011101111110111110011;
            'd127: data <= 32'b01101011011011011011111111010010;
            'd128: data <= 32'b00111010010011001000000111001101;
            'd129: data <= 32'b10010001000101000001100000001100;
            'd130: data <= 32'b00010001001101010010011000010011;
            'd131: data <= 32'b01000001001011111100001111101100;
            'd132: data <= 32'b01001111111000011011111001011111;
            'd133: data <= 32'b01100111101000100011010110010111;
            'd134: data <= 32'b11011100110011001000100001000100;
            'd135: data <= 32'b11101010001110010010111000010111;
            'd136: data <= 32'b10010111010101111001001111000100;
            'd137: data <= 32'b11110010111100100101010110100111;
            'd138: data <= 32'b11001111100000101111110001111110;
            'd139: data <= 32'b11001110010001110111101000111101;
            'd140: data <= 32'b11110000101011001100100001100100;
            'd141: data <= 32'b10110100111001111011101001011101;
            'd142: data <= 32'b11100110001010110011001000011001;
            'd143: data <= 32'b01110011100101011110011001110011;
            'd144: data <= 32'b10010110101000001100000001100000;
            'd145: data <= 32'b10101100100110000001100110000001;
            'd146: data <= 32'b01110100110100011001111001001111;
            'd147: data <= 32'b00100010011111111010001111011100;
            'd148: data <= 32'b11100111011001100100010000100010;
            'd149: data <= 32'b10101101011111100101010000101010;
            'd150: data <= 32'b00110101101010110011101110010000;
            'd151: data <= 32'b10000101100000110000101110001000;
            'd152: data <= 32'b11100010110010101000110001000110;
            'd153: data <= 32'b11111001001010011100011111101110;
            'd154: data <= 32'b00110111110100110110101110111000;
            'd155: data <= 32'b11101000001111000010100000010100;
            'd156: data <= 32'b00011100011110011010011111011110;
            'd157: data <= 32'b01110101111000101011110001011110;
            'd158: data <= 32'b11011111000111010001011000001011;
            'd159: data <= 32'b01101110011101101010110111011011;
            'd160: data <= 32'b01000111001110111101101111100000;
            'd161: data <= 32'b11110001010101100110010000110010;
            'd162: data <= 32'b00011010010011100111010000111010;
            'd163: data <= 32'b01110001000111100001010000001010;
            'd164: data <= 32'b00011101110110111001001001001001;
            'd165: data <= 32'b00101001000010100000110000000110;
            'd166: data <= 32'b11000101011011000100100000100100;
            'd167: data <= 32'b10001001111001001011100001011100;
            'd168: data <= 32'b01101111010111011001111111000010;
            'd169: data <= 32'b10110111011011101011110111010011;
            'd170: data <= 32'b01100010111011110100001110101100;
            'd171: data <= 32'b00001110101001101100010001100010;
            'd172: data <= 32'b10101010101010000011100110010001;
            'd173: data <= 32'b00011000101001000011000110010101;
            'd174: data <= 32'b10111110001101111101001111100100;
            'd175: data <= 32'b00011011100010111111001001111001;
            'd176: data <= 32'b11111100001100101101010111100111;
            'd177: data <= 32'b01010110010000111000101111001000;
            'd178: data <= 32'b00111110010110010110111000110111;
            'd179: data <= 32'b01001011101101111101101001101101;
            'd180: data <= 32'b11000110100011000000000110001101;
            'd181: data <= 32'b11010010011001001011000111010101;
            'd182: data <= 32'b01111001110100101001110001001110;
            'd183: data <= 32'b00100000111000000100100110101001;
            'd184: data <= 32'b10011010101101001101100001101100;
            'd185: data <= 32'b11011011111110101010110001010110;
            'd186: data <= 32'b11000000000001111111001111110100;
            'd187: data <= 32'b11111110001001011100111111101010;
            'd188: data <= 32'b01111000101011111100101001100101;
            'd189: data <= 32'b11001101100011101111010001111010;
            'd190: data <= 32'b01011010111010010100011110101110;
            'd191: data <= 32'b11110100000110000001000000001000;
            'd192: data <= 32'b00011111110101010110111110111010;
            'd193: data <= 32'b11011101100010001111000001111000;
            'd194: data <= 32'b10101000011011110100101000100101;
            'd195: data <= 32'b00110011011100100101110000101110;
            'd196: data <= 32'b10001000001001000011100000011100;
            'd197: data <= 32'b00000111111100010101011110100110;
            'd198: data <= 32'b11000111110001110111001110110100;
            'd199: data <= 32'b00110001010100011001011111000110;
            'd200: data <= 32'b10110001001000111100101111101000;
            'd201: data <= 32'b00010010011111001010000111011101;
            'd202: data <= 32'b00010000100111001110100001110100;
            'd203: data <= 32'b01011001001000010011111000011111;
            'd204: data <= 32'b00100111110111011001011001001011;
            'd205: data <= 32'b10000000110111000110000110111101;
            'd206: data <= 32'b11101100100001100000110110001011;
            'd207: data <= 32'b01011111100001010000111110001010;
            'd208: data <= 32'b01100000100100001110000001110000;
            'd209: data <= 32'b01010001010000100111110000111110;
            'd210: data <= 32'b01111111110001000111000110110101;
            'd211: data <= 32'b10101001101010101100110001100110;
            'd212: data <= 32'b00011001110110001001000001001000;
            'd213: data <= 32'b10110101000001010000011000000011;
            'd214: data <= 32'b01001010000000011111011111110110;
            'd215: data <= 32'b00001101000100100001110000001110;
            'd216: data <= 32'b00101101101000111100001001100001;
            'd217: data <= 32'b11100101010111110110101000110101;
            'd218: data <= 32'b01111010111110011010111001010111;
            'd219: data <= 32'b10011111110100000110100110111001;
            'd220: data <= 32'b10010011100100010001011110000110;
            'd221: data <= 32'b11001001010110001001100111000001;
            'd222: data <= 32'b10011100001001110011101000011101;
            'd223: data <= 32'b11101111101110010010011110011110;
            'd224: data <= 32'b10100000001110001101100111100001;
            'd225: data <= 32'b11100000000100111110101111111000;
            'd226: data <= 32'b00111011101100110010101110011000;
            'd227: data <= 32'b01001101001100110010001000010001;
            'd228: data <= 32'b10101110101110111101001001101001;
            'd229: data <= 32'b00101010011100001010100111011001;
            'd230: data <= 32'b11110101100010010000011110001110;
            'd231: data <= 32'b10110000101001110011001110010100;
            'd232: data <= 32'b11001000101101100010110110011011;
            'd233: data <= 32'b11101011001000100011110000011110;
            'd234: data <= 32'b10111011100100100001010110000111;
            'd235: data <= 32'b00111100001000001100100111101001;
            'd236: data <= 32'b10000011010010011000011111001110;
            'd237: data <= 32'b01010011111111111010101001010101;
            'd238: data <= 32'b10011001011110000101000000101000;
            'd239: data <= 32'b01100001011110101010010111011111;
            'd240: data <= 32'b00010111100011110000001110001100;
            'd241: data <= 32'b00101011111110000101100110100001;
            'd242: data <= 32'b00000100100000000000100110001001;
            'd243: data <= 32'b01111110000101110001101000001101;
            'd244: data <= 32'b10111010110110100110010110111111;
            'd245: data <= 32'b01110111001100011101011111100110;
            'd246: data <= 32'b11010110110001101000010001000010;
            'd247: data <= 32'b00100110101110001101000001101000;
            'd248: data <= 32'b11100001110000111000001001000001;
            'd249: data <= 32'b01101001101100000010100110011001;
            'd250: data <= 32'b00010100011101110101101000101101;
            'd251: data <= 32'b01100011000100010001111000001111;
            'd252: data <= 32'b01010101110010110111101110110000;
            'd253: data <= 32'b00100001111111001010100001010100;
            'd254: data <= 32'b00001100110101100110110110111011;
            'd255: data <= 32'b01111101001110100010110000010110;
            'd256: data <= 32'b01010000101001111111010001010001;
            'd257: data <= 32'b01010011011001010100000101111110;
            'd258: data <= 32'b11000011101001000001011100011010;
            'd259: data <= 32'b10010110010111100010011100111010;
            'd260: data <= 32'b11001011011010111010101100111011;
            'd261: data <= 32'b11110001010001011001110100011111;
            'd262: data <= 32'b10101011010110001111101010101100;
            'd263: data <= 32'b10010011000000111110001101001011;
            'd264: data <= 32'b01010101111110100011000000100000;
            'd265: data <= 32'b11110110011011010111011010101101;
            'd266: data <= 32'b10010001011101101100110010001000;
            'd267: data <= 32'b00100101010011000000001011110101;
            'd268: data <= 32'b11111100110101111110010101001111;
            'd269: data <= 32'b11010111110010110010101011000101;
            'd270: data <= 32'b10000000010001000011010100100110;
            'd271: data <= 32'b10001111101000110110001010110101;
            'd272: data <= 32'b01001001010110101011000111011110;
            'd273: data <= 32'b01100111000110111011101000100101;
            'd274: data <= 32'b10011000000011101110101001000101;
            'd275: data <= 32'b11100001110000001111111001011101;
            'd276: data <= 32'b00000010011101010010111111000011;
            'd277: data <= 32'b00010010111100000100110010000001;
            'd278: data <= 32'b10100011100101110100011010001101;
            'd279: data <= 32'b11000110111110011101001101101011;
            'd280: data <= 32'b11100111010111111000111100000011;
            'd281: data <= 32'b10010101100111001001001000010101;
            'd282: data <= 32'b11101011011110100110110110111111;
            'd283: data <= 32'b11011010010110010101001010010101;
            'd284: data <= 32'b00101101100000111011111011010100;
            'd285: data <= 32'b11010011001000010111010001011000;
            'd286: data <= 32'b00101001011010011110000001001001;
            'd287: data <= 32'b01000100110010001100100110001110;
            'd288: data <= 32'b01101010100010011100001001110101;
            'd289: data <= 32'b01111000011110011000111011110100;
            'd290: data <= 32'b01101011001111100101100010011001;
            'd291: data <= 32'b11011101011100011011100100100111;
            'd292: data <= 32'b10110110010011111110000110111110;
            'd293: data <= 32'b00010111101011011000100011110000;
            'd294: data <= 32'b01100110101011000010000011001001;
            'd295: data <= 32'b10110100001110101100111001111101;
            'd296: data <= 32'b00011000010010101101111101100011;
            'd297: data <= 32'b10000010001100010001101011100101;
            'd298: data <= 32'b01100000001100110101000110010111;
            'd299: data <= 32'b01000101011111110101001101100010;
            'd300: data <= 32'b11100000011101110110010010110001;
            'd301: data <= 32'b10000100101011100110101110111011;
            'd302: data <= 32'b00011100101000001000000111111110;
            'd303: data <= 32'b10010100001010110000100011111001;
            'd304: data <= 32'b01011000011010000100100001110000;
            'd305: data <= 32'b00011001111111010100010110001111;
            'd306: data <= 32'b10000111011011001101111010010100;
            'd307: data <= 32'b10110111111110000111101101010010;
            'd308: data <= 32'b00100011110100110111001110101011;
            'd309: data <= 32'b11100010000000100100101101110010;
            'd310: data <= 32'b01010111100011110001111111100011;
            'd311: data <= 32'b00101010101010110101010101100110;
            'd312: data <= 32'b00000111001010001110101110110010;
            'd313: data <= 32'b00000011110000101011010100101111;
            'd314: data <= 32'b10011010011110111100010110000110;
            'd315: data <= 32'b10100101000010000011011111010011;
            'd316: data <= 32'b11110010100001110010100000110000;
            'd317: data <= 32'b10110010101001011011111100100011;
            'd318: data <= 32'b10111010011010100000001100000010;
            'd319: data <= 32'b01011100100000100001011011101101;
            'd320: data <= 32'b00101011000111001100111110001010;
            'd321: data <= 32'b10010010101101000111100110100111;
            'd322: data <= 32'b11110000111100100000011111110011;
            'd323: data <= 32'b10100001111000100110100101001110;
            'd324: data <= 32'b11001101111101001101101001100101;
            'd325: data <= 32'b11010101101111100000010100000110;
            'd326: data <= 32'b00011111011000100011010011010001;
            'd327: data <= 32'b10001010111111101010011011000100;
            'd328: data <= 32'b10011101010100110010111000110100;
            'd329: data <= 32'b10100000010101011111001110100010;
            'd330: data <= 32'b00110010111000011000101000000101;
            'd331: data <= 32'b01110101111010111111011010100100;
            'd332: data <= 32'b00111001111011001000001100001011;
            'd333: data <= 32'b10101010111011110110000001000000;
            'd334: data <= 32'b00000110100111110111000101011110;
            'd335: data <= 32'b01010001000100000110111010111101;
            'd336: data <= 32'b11111001100010100010000100111110;
            'd337: data <= 32'b00111101000001101101110110010110;
            'd338: data <= 32'b10101110000001010011111011011101;
            'd339: data <= 32'b01000110101111011110011001001101;
            'd340: data <= 32'b10110101100011010101010010010001;
            'd341: data <= 32'b00000101010111011100010001110001;
            'd342: data <= 32'b01101111110101000000011000000100;
            'd343: data <= 32'b11111111000101010101000001100000;
            'd344: data <= 32'b00100100111110111001100000011001;
            'd345: data <= 32'b10010111111010011011110111010110;
            'd346: data <= 32'b11001100010000110100000010001001;
            'd347: data <= 32'b01110111100111101101100101100111;
            'd348: data <= 32'b10111101010000101110100010110000;
            'd349: data <= 32'b10001000100010111000100100000111;
            'd350: data <= 32'b00111000010110110001100111100111;
            'd351: data <= 32'b11011011111011101100100001111001;
            'd352: data <= 32'b01000111000010100111110010100001;
            'd353: data <= 32'b11101001000011110100001001111100;
            'd354: data <= 32'b11001001000111101000010011111000;
            'd355: data <= 32'b00000000000000000000000000000000;
            'd356: data <= 32'b10000011100001101000000000001001;
            'd357: data <= 32'b01001000111011010010101100110010;
            'd358: data <= 32'b10101100011100000001000100011110;
            'd359: data <= 32'b01001110011100100101101001101100;
            'd360: data <= 32'b11111011111111110000111011111101;
            'd361: data <= 32'b01010110001110001000010100001111;
            'd362: data <= 32'b00011110110101011010111000111101;
            'd363: data <= 32'b00100111001110010010110100110110;
            'd364: data <= 32'b01100100110110010000111100001010;
            'd365: data <= 32'b00100001101001100101110001101000;
            'd366: data <= 32'b11010001010101000101101110011011;
            'd367: data <= 32'b00111010001011100011011000100100;
            'd368: data <= 32'b10110001011001110000101000001100;
            'd369: data <= 32'b00001111111001110101011110010011;
            'd370: data <= 32'b11010010100101101110111010110100;
            'd371: data <= 32'b10011110100100011001101100011011;
            'd372: data <= 32'b01001111110001011100000010000000;
            'd373: data <= 32'b10100010001000001101110001100001;
            'd374: data <= 32'b01101001010010110111011101011010;
            'd375: data <= 32'b00010110000110100001001000011100;
            'd376: data <= 32'b00001010101110101001001111100010;
            'd377: data <= 32'b11100101001010101010000011000000;
            'd378: data <= 32'b01000011111000000010001000111100;
            'd379: data <= 32'b00011101000101110001101100010010;
            'd380: data <= 32'b00001011000011010000100100001110;
            'd381: data <= 32'b10101101110001111000101111110010;
            'd382: data <= 32'b10111001101010001011011000101101;
            'd383: data <= 32'b11001000101010010001111000010100;
            'd384: data <= 32'b10000101000110011111000101010111;
            'd385: data <= 32'b01001100000001110111010110101111;
            'd386: data <= 32'b10111011110111011001100111101110;
            'd387: data <= 32'b11111101011000000111111110100011;
            'd388: data <= 32'b10011111001001100000000111110111;
            'd389: data <= 32'b10111100111101010111001001011100;
            'd390: data <= 32'b11000101001110110110011001000100;
            'd391: data <= 32'b00110100011111101111101101011011;
            'd392: data <= 32'b01110110001010010100001110001011;
            'd393: data <= 32'b11011100110001100010001111001011;
            'd394: data <= 32'b01101000111111001110110110110110;
            'd395: data <= 32'b01100011111100011110010010111000;
            'd396: data <= 32'b11001010110111000011000111010111;
            'd397: data <= 32'b00010000100001010110001101000010;
            'd398: data <= 32'b01000000001000101001011100010011;
            'd399: data <= 32'b00100000000100011100011010000100;
            'd400: data <= 32'b01111101001001000100101010000101;
            'd401: data <= 32'b11111000001111011011101111010010;
            'd402: data <= 32'b00010001001100101111100110101110;
            'd403: data <= 32'b01101101101000010010100111000111;
            'd404: data <= 32'b01001011001011111001111000011101;
            'd405: data <= 32'b11110011001100001011001011011100;
            'd406: data <= 32'b11101100010100101000011000001101;
            'd407: data <= 32'b11010000111000111100000101110111;
            'd408: data <= 32'b01101100000101101011001100101011;
            'd409: data <= 32'b10011001101110010111000010101001;
            'd410: data <= 32'b11111010010010001001010000010001;
            'd411: data <= 32'b00100010011001001110100101000111;
            'd412: data <= 32'b11000100100011001111110010101000;
            'd413: data <= 32'b00011010001111111111000010100000;
            'd414: data <= 32'b11011000001011000111110101010110;
            'd415: data <= 32'b11101111100100000011001100100010;
            'd416: data <= 32'b11000111010011100100100110000111;
            'd417: data <= 32'b11000001110100010011100011011001;
            'd418: data <= 32'b11111110101000101100101010001100;
            'd419: data <= 32'b00110110000010111101010010011000;
            'd420: data <= 32'b11001111100000011111010110100110;
            'd421: data <= 32'b00101000110111100111101010100101;
            'd422: data <= 32'b00100110100011101011011111011010;
            'd423: data <= 32'b10100100101111111010110100111111;
            'd424: data <= 32'b11100100100111010011101000101100;
            'd425: data <= 32'b00001101100100100111100001010000;
            'd426: data <= 32'b10011011110011000101111101101010;
            'd427: data <= 32'b01100010010001100111111001010100;
            'd428: data <= 32'b11000010000100111000110111110110;
            'd429: data <= 32'b11101000101110001101100010010000;
            'd430: data <= 32'b01011110111101110011100100101110;
            'd431: data <= 32'b11110101101011111100001110000010;
            'd432: data <= 32'b10111110100000000101110110011111;
            'd433: data <= 32'b01111100100100111101000001101001;
            'd434: data <= 32'b10101001001011011101010101101111;
            'd435: data <= 32'b10110011000100100010010111001111;
            'd436: data <= 32'b00111011100110011010110011001000;
            'd437: data <= 32'b10100111011111010001100000010000;
            'd438: data <= 32'b01101110011000111001110011101000;
            'd439: data <= 32'b01111011101110110011101111011011;
            'd440: data <= 32'b00001001011110000010011011001101;
            'd441: data <= 32'b11110100000110000101100101101110;
            'd442: data <= 32'b00000001101101111001101011101100;
            'd443: data <= 32'b10101000100110100100111110000011;
            'd444: data <= 32'b01100101011011101001010111100110;
            'd445: data <= 32'b01111110111001101111111110101010;
            'd446: data <= 32'b00001000110011111011110000100001;
            'd447: data <= 32'b11100110111010000001010111101111;
            'd448: data <= 32'b11011001100110111110011110111010;
            'd449: data <= 32'b11001110001101100110111101001010;
            'd450: data <= 32'b11010100000010011001111111101010;
            'd451: data <= 32'b11010110011111001011000000101001;
            'd452: data <= 32'b10101111101100101010010000110001;
            'd453: data <= 32'b00110001001000110011111100101010;
            'd454: data <= 32'b00110000100101001010010111000110;
            'd455: data <= 32'b11000000011001101010001000110101;
            'd456: data <= 32'b00110111101111000100111001110100;
            'd457: data <= 32'b10100110110010101000001011111100;
            'd458: data <= 32'b10110000110100001001000011100000;
            'd459: data <= 32'b00010101110110001010011100110011;
            'd460: data <= 32'b01001010100110000000010011110001;
            'd461: data <= 32'b11110111110110101110110001000001;
            'd462: data <= 32'b00001110010100001100110101111111;
            'd463: data <= 32'b00101111111101101001000100010111;
            'd464: data <= 32'b10001101110101100100110101110110;
            'd465: data <= 32'b01001101101100001110111101000011;
            'd466: data <= 32'b01010100010011011010101011001100;
            'd467: data <= 32'b11011111000001001001011011100100;
            'd468: data <= 32'b11100011101101011101000110011110;
            'd469: data <= 32'b00011011100010000110101001001100;
            'd470: data <= 32'b10111000000111110010110011000001;
            'd471: data <= 32'b01111111010100010110010101000110;
            'd472: data <= 32'b00000100111010100101111010011101;
            'd473: data <= 32'b01011101001101011000110000000001;
            'd474: data <= 32'b01110011011101001000011111111010;
            'd475: data <= 32'b00101110010000010000101111111011;
            'd476: data <= 32'b01011010000111010110011110110011;
            'd477: data <= 32'b01010010110100101101101110010010;
            'd478: data <= 32'b00110011010101100001000011101001;
            'd479: data <= 32'b00010011010001111101011001101101;
            'd480: data <= 32'b10001100011000011101011110011010;
            'd481: data <= 32'b01111010000011001010000100110111;
            'd482: data <= 32'b10001110000101001111100001011001;
            'd483: data <= 32'b10001001001111000001001111101011;
            'd484: data <= 32'b11101110001001111010100111001110;
            'd485: data <= 32'b00110101110010010110000110110111;
            'd486: data <= 32'b11101101111001010001110011100001;
            'd487: data <= 32'b00111100101100010100011101111010;
            'd488: data <= 32'b01011001110111111101001010011100;
            'd489: data <= 32'b00111111011100111111001001010101;
            'd490: data <= 32'b01111001110011100001010000011000;
            'd491: data <= 32'b10111111001101111100011101110011;
            'd492: data <= 32'b11101010110011011111011101010011;
            'd493: data <= 32'b01011011101010101111110101011111;
            'd494: data <= 32'b00010100011011110011110111011111;
            'd495: data <= 32'b10000110110110110100010001111000;
            'd496: data <= 32'b10000001111100111010111111001010;
            'd497: data <= 32'b00111110110001000110100010111001;
            'd498: data <= 32'b00101100001101000010010000111000;
            'd499: data <= 32'b01011111010000001010001111000010;
            'd500: data <= 32'b01110010110000110001110100010110;
            'd501: data <= 32'b00001100001001011110001010111100;
            'd502: data <= 32'b10001011010010010011110000101000;
            'd503: data <= 32'b01000001100101010000110111111111;
            'd504: data <= 32'b01110001000000011010100000111001;
            'd505: data <= 32'b11011110101100110000110000001000;
            'd506: data <= 32'b10011100111001001011010011011000;
            'd507: data <= 32'b10010000110000010101011001100100;
            'd508: data <= 32'b01100001100001001100101101111011;
            'd509: data <= 32'b01110000101101100011001011010101;
            'd510: data <= 32'b01110100010111000110110001001000;
            'd511: data <= 32'b01000010010101111011100011010000;


            default: data <= 32'h0;
        endcase
    end else begin
        data <= data;
    end
end

endmodule
`resetall
