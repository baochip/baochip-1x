// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: SHL-0.51
//
// This file has been modified by CrossBar, Inc.

// Copyright 2015-2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

`undef SPI_STD          
`undef SPI_QUAD_TX      
`undef SPI_QUAD_RX      
`undef SPI_CMD_CFG      
`undef SPI_CMD_SOT      
`undef SPI_CMD_SEND_CMD 
`undef SPI_CMD_DUMMY    
`undef SPI_CMD_WAIT     
`undef SPI_CMD_TX_DATA  
`undef SPI_CMD_RX_DATA  
`undef SPI_CMD_RPT      
`undef SPI_CMD_EOT      
`undef SPI_CMD_RPT_END  
`undef SPI_CMD_RX_CHECK 
`undef SPI_CMD_FULL_DUPL
`undef SPI_CMD_SETUP_UCA
`undef SPI_CMD_SETUP_UCS
`undef REG_RX_SADDR     
`undef REG_RX_SIZE      
`undef REG_RX_CFG       
`undef REG_RX_INTCFG    
`undef REG_TX_SADDR     
`undef REG_TX_SIZE      
`undef REG_TX_CFG       
`undef REG_TX_INTCFG    
`undef REG_CMD_SADDR    
`undef REG_CMD_SIZE     
`undef REG_CMD_CFG      
`undef REG_CMD_INTCFG   
`undef REG_STATUS       
`undef SPI_WAIT_EVT     
`undef SPI_WAIT_CYC     
`undef SPI_WAIT_GP      