// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

//`include "ips/nic400_1/logical/nic400_1/amib_m0/verilog/nic400_amib_m0_defs_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m0/verilog/nic400_amib_m0_undefs_1.v"
`include "ips/nic400_1/logical/nic400_1/amib_m0/verilog/nic400_amib_m0_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m0/verilog/Ahb.v"
////`include "ips/nic400_1/logical/nic400_1/amib_m0/verilog/Ahb_undefs.v"
`include "ips/nic400_1/logical/nic400_1/amib_m0/verilog/nic400_amib_m0_chan_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/amib_m1/verilog/nic400_amib_m1_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m1/verilog/nic400_amib_m1_defs_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m1/verilog/nic400_amib_m1_undefs_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m1/verilog/Ahb.v"
`include "ips/nic400_1/logical/nic400_1/amib_m1/verilog/nic400_amib_m1_chan_slice_1.v"
////`include "ips/nic400_1/logical/nic400_1/amib_m1/verilog/Ahb_undefs.v"
`include "ips/nic400_1/logical/nic400_1/amib_m2/verilog/nic400_amib_m2_chan_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m2/verilog/nic400_amib_m2_undefs_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m2/verilog/Ahb.v"
`include "ips/nic400_1/logical/nic400_1/amib_m2/verilog/nic400_amib_m2_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m2/verilog/nic400_amib_m2_defs_1.v"
////`include "ips/nic400_1/logical/nic400_1/amib_m2/verilog/Ahb_undefs.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m3/verilog/nic400_amib_m3_defs_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m3/verilog/nic400_amib_m3_undefs_1.v"
`include "ips/nic400_1/logical/nic400_1/amib_m3/verilog/nic400_amib_m3_chan_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/amib_m3/verilog/Ahb.v"
////`include "ips/nic400_1/logical/nic400_1/amib_m3/verilog/Ahb_undefs.v"
`include "ips/nic400_1/logical/nic400_1/amib_m3/verilog/nic400_amib_m3_1.v"

`include "ips/nic400_1/logical/nic400_1/asib_s0/verilog/nic400_asib_s0_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s0/verilog/nic400_asib_s0_maskcntl_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s0/verilog/nic400_asib_s0_chan_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s0/verilog/nic400_asib_s0_rd_ss_cdas_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s0/verilog/nic400_asib_s0_wr_ss_cdas_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s0/verilog/nic400_asib_s0_decode_1.v"

`include "ips/nic400_1/logical/nic400_1/asib_s2/verilog/nic400_asib_s2_rd_ss_cdas_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s2/verilog/nic400_asib_s2_decode_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s2/verilog/nic400_asib_s2_wr_ss_cdas_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s2/verilog/nic400_asib_s2_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s2/verilog/nic400_asib_s2_chan_slice_1.v"

`include "ips/nic400_1/logical/nic400_1/asib_s3/verilog/nic400_asib_s3_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s3/verilog/nic400_asib_s3_maskcntl_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s3/verilog/nic400_asib_s3_chan_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s3/verilog/nic400_asib_s3_rd_ss_cdas_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s3/verilog/nic400_asib_s3_wr_ss_cdas_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s3/verilog/nic400_asib_s3_decode_1.v"

`include "ips/nic400_1/logical/nic400_1/asib_s4/verilog/nic400_asib_s4_rd_ss_cdas_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s4/verilog/nic400_asib_s4_decode_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s4/verilog/nic400_asib_s4_wr_ss_cdas_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s4/verilog/nic400_asib_s4_1.v"
`include "ips/nic400_1/logical/nic400_1/asib_s4/verilog/nic400_asib_s4_chan_slice_1.v"







//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_2_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_blayer_1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml4_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml4_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_map_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml3_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml4_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_blayer_0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_st_tt_s0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_2_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml2_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml3_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_ss_tt_s1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_3_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_3_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_4_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_ss_tt_s1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml3_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml2_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml2_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_lrg_arb_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml3_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_build_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_ss_tt_s0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml2_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml4_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml1_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml2_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml3_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_qv_cmp_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_0_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml4_1.v"
//`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_1_1.v"


`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_arb_ml4_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml4_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_lrg_arb_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml4_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_blayer_0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_blayer_1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_blayer_2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_blayer_3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_build_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_map_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_4_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_qv_cmp_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_ss_tt_s0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_ss_tt_s1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_ss_tt_s2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_ss_tt_s3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml4_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml2_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml4_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_ss_tt_s1_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_ss_tt_s3_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_st_tt_s0_1.v"
`include "ips/nic400_1/logical/nic400_1/busmatrix_bm0/verilog/nic400_bm0_wr_st_tt_s2_1.v"



//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_launch_data_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_sync_flop_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_corrupt_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_capt_nosync_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_reset_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_comb_and2_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_random_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_comb_or2_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_syncn_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_bypass_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_capt_sync_1.v"
`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_comb_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_launch_gry_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_corrupt_gry_1.v"
//`include "ips/nic400_1/logical/nic400_1/cdc_blocks/verilog/nic400_cdc_comb_or3_1.v"
//`include "ips/nic400_1/logical/nic400_1/default_slave_ds_1/verilog/nic400_default_slave_ds_1_undefs_1.v"
//`include "ips/nic400_1/logical/nic400_1/default_slave_ds_1/verilog/nic400_default_slave_ds_1_defs_1.v"
`include "ips/nic400_1/logical/nic400_1/default_slave_ds_1/verilog/nic400_default_slave_ds_1_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_slave_domain_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_b_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_chan_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_w_fifo_wr_mux2_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_ar_fifo_wr_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_r_fifo_wr_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_b_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_undefs_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_upsize_wr_resp_block_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_upsize_resp_cam_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_aw_fifo_wr_mux_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_w_fifo_wr_mux_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_w_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_aw_fifo_fn_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_maskcntl_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_b_fifo_wr_mux2_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_aw_fifo_wr_mux2_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_upsize_rd_cam_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_w_fifo_sync_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_ar_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_ar_fifo_fn_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_w_fifo_wr_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_ar_fifo_sync_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_aw_fifo_rd_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_upsize_rd_addr_fmt_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_b_fifo_wr_mux_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_r_fifo_wr_mux_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_aw_fifo_sync_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_upsize_wr_cntrl_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_b_fifo_wr_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_r_fifo_wr_mux2_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_ar_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_defs_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_b_fifo_fn_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_r_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_r_fifo_fn_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_w_fifo_fn_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_upsize_rd_chan_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_upsize_wr_merge_buffer_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_upsize_wr_addr_fmt_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_ar_fifo_wr_mux2_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_r_fifo_sync_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_master_domain_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s2_ib/verilog/nic400_ib_s2_ib_aw_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/verilog/Axi4PC/Axi4PC_undefs.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/verilog/Axi4PC/Axi4PC_message_undefs.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/verilog/Axi4PC/Axi4PC_no_coverage_macros.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/verilog/Axi4PC/Axi4PC_defs.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/verilog/Axi4PC/Axi4PC_coverage_undefs.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/verilog/Axi4PC/Axi4PC_message_defs.v"
`include "ips/nic400_1/logical/nic400_1/nic400/verilog/nic400_1.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/verilog/Axi/Axi.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/verilog/Axi/Axi_undefs.v"
`include "ips/nic400_1/logical/nic400_1/nic400/verilog/nic400_cd_clk1_1.v"
`include "ips/nic400_1/logical/nic400_1/nic400/verilog/nic400_cd_clk0_1.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/validation/shared/tbench/tbench.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/validation/shared/tb_components/clk_reset_if.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/validation/shared/tb_components/config_if.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/validation/shared/tb_components/ahb_aux.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/validation/shared/tb_components/FrmEventDistributor.v"
//`include "ips/nic400_1/logical/nic400_1/nic400/validation/shared/tb_components/apb_aux.v"
`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_rev_regd_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_fwd_regd_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_ful_regd_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/reg_slice_axi_undefs.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_wr4_reg_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_buf_reg_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_ax_reg_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_wr_reg_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_ax4_reg_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_reg_slice_axi_1.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/reg_slice_axi_defs.v"
//`include "ips/nic400_1/logical/nic400_1/reg_slice/verilog/nic400_rd_reg_slice_1.v"

//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_slave_domain_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_b_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_w_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_ar_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_r_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_b_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_upsize_wr_resp_block_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_upsize_resp_cam_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_aw_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_w_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_w_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_maskcntl_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_b_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_aw_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_upsize_rd_cam_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_w_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_ar_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_w_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_ar_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_aw_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_upsize_rd_addr_fmt_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_b_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_r_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_aw_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_upsize_wr_cntrl_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_b_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_r_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_ar_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_r_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_upsize_rd_chan_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_upsize_wr_merge_buffer_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_upsize_wr_addr_fmt_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_ar_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_r_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_master_domain_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s3_ib/verilog/nic400_ib_s3_ib_aw_fifo_wr_1.v"

//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_chan_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_maskcntl_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_master_domain_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_slave_domain_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_addr_fmt_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_cam_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_chan_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_resp_cam_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_addr_fmt_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_cntrl_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_merge_buffer_1.v"


`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_chan_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_maskcntl_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_master_domain_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_slave_domain_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_addr_fmt_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_cam_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_chan_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_resp_cam_slice_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_addr_fmt_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_cntrl_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_merge_buffer_1.v"
`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_resp_block_1.v"


//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_slave_domain_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_b_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_w_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_ar_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_r_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_b_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_resp_block_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_resp_cam_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_aw_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_w_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_w_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_maskcntl_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_b_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_aw_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_cam_slice_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_w_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_ar_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_w_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_ar_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_aw_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_addr_fmt_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_b_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_r_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_aw_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_cntrl_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_b_fifo_wr_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_r_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_ar_fifo_wr_mux_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_r_fifo_rd_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_rd_chan_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_merge_buffer_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_upsize_wr_addr_fmt_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_ar_fifo_wr_mux2_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_r_fifo_sync_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_master_domain_1.v"
//`include "ips/nic400_1/logical/nic400_1/ib_s4_ib/verilog/nic400_ib_s4_ib_aw_fifo_wr_1.v"