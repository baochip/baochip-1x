// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

// -----------------------------------------------------------------------------
// Auto-Generated by:        __   _ __      _  __
//                          / /  (_) /____ | |/_/
//                         / /__/ / __/ -_)>  <
//                        /____/_/\__/\__/_/|_|
//                     Build your hardware, easily!
//                   https://github.com/enjoy-digital/litex
//
// Filename   : cdc_blinded.v
// Device     : generic
// LiteX sha1 : 37d630db
// Date       : 2023-05-10 14:56:55
//------------------------------------------------------------------------------

`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// Module
//------------------------------------------------------------------------------

module cdc_blinded (
    input  wire          reset,
    input  wire          clk_a,
    input  wire          clk_b,
    input  wire          in_a,
    output wire          out_b
);


//------------------------------------------------------------------------------
// Signals
//------------------------------------------------------------------------------

wire          a_clk;
wire          a_rst;
wire          b_clk;
wire          b_rst;
wire          i;
wire          o;
wire          ps_i;
wire          ps_o;
reg           ps_toggle_i;
wire          ps_toggle_o;
reg           ps_toggle_o_r;
wire          ps_ack_i;
wire          ps_ack_o;
reg           ps_ack_toggle_i;
wire          ps_ack_toggle_o;
reg           ps_ack_toggle_o_r;
reg           blind;
reg           multiregimpl00;
reg           multiregimpl01;
reg           multiregimpl10;
reg           multiregimpl11;

//------------------------------------------------------------------------------
// Combinatorial Logic
//------------------------------------------------------------------------------

assign a_clk = clk_a;
assign a_rst = reset;
assign b_clk = clk_b;
assign b_rst = reset;
assign i = in_a;
assign out_b = o;
assign ps_i = (i & (~blind));
assign ps_ack_i = ps_o;
assign o = ps_o;
assign ps_o = (ps_toggle_o ^ ps_toggle_o_r);
assign ps_ack_o = (ps_ack_toggle_o ^ ps_ack_toggle_o_r);
assign ps_toggle_o = multiregimpl01;
assign ps_ack_toggle_o = multiregimpl11;


//------------------------------------------------------------------------------
// Synchronous Logic
//------------------------------------------------------------------------------

always @(posedge a_clk) begin
    if (i) begin
        blind <= 1'd1;
    end
    if (ps_ack_o) begin
        blind <= 1'd0;
    end
    if (a_rst) begin
        ps_toggle_i <= 0;
    end else if (ps_i) begin
        ps_toggle_i <= (~ps_toggle_i);
    end
    ps_ack_toggle_o_r <= ps_ack_toggle_o;
    if (a_rst) begin
        blind <= 1'd0;
    end
    multiregimpl10 <= ps_ack_toggle_i;
    multiregimpl11 <= multiregimpl10;
end

always @(posedge b_clk) begin
    ps_toggle_o_r <= ps_toggle_o;
    if (b_rst) begin
        ps_ack_toggle_i <= 0;
    end else if (ps_ack_i) begin
        ps_ack_toggle_i <= (~ps_ack_toggle_i);
    end
    multiregimpl00 <= ps_toggle_i;
    multiregimpl01 <= multiregimpl00;
end


//------------------------------------------------------------------------------
// Specialized Logic
//------------------------------------------------------------------------------

endmodule

// -----------------------------------------------------------------------------
//  Auto-Generated by LiteX on 2023-05-10 14:56:55.
//------------------------------------------------------------------------------
