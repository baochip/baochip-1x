// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

`include "template.sv"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml1_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_wr_st_tt_s0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_add_sel_ml1_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_rd_st_tt_s0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_ml_map_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml1_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_ml_build_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_1_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_rd_wr_arb_0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_maskcntl_ml0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_ml_blayer_0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_ret_sel_ml0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_wr_sel_ml1_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/busmatrix_bm0/verilog/nic400_bm0_ml_mlayer_0_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/default_slave_ds_1/verilog/nic400_default_slave_ds_1_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/default_slave_ds_1/verilog/nic400_default_slave_ds_1_undefs_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/default_slave_ds_1/verilog/nic400_default_slave_ds_1_defs_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Axi4PC/Axi4PC_undefs.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Axi4PC/Axi4PC_message_undefs.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Axi4PC/Axi4PC_no_coverage_macros.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Axi4PC/Axi4PC_defs.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Axi4PC/Axi4PC_coverage_undefs.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Axi4PC/Axi4PC_message_defs.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/AhbPC/AhbPC.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Axi/Axi.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Axi/Axi_undefs.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Ahb/AhbDefns.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/Ahb/AhbDefns_undefs.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/nic400/verilog/nic400_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_fwd_regd_slice_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_ax4_reg_slice_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_rev_regd_slice_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_ax_reg_slice_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_wr4_reg_slice_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/reg_slice_axi_undefs.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_buf_reg_slice_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_wr_reg_slice_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_rd_reg_slice_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_ful_regd_slice_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/reg_slice_axi_defs.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/reg_slice/verilog/nic400_reg_slice_axi_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_comb_mux2_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_corrupt_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_comb_or3_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_launch_gry_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_corrupt_gry_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_launch_data_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_bypass_sync_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_comb_or2_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_capt_sync_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_random_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_comb_and2_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_reset_sync_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_cdc_capt_nosync_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_sync_flop_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/cdc_blocks/verilog/nic400_syncn_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_ahb_undefs_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_defs_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_undefs_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_ahb_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_chan_slice_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_itb_to_axi_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_rd_ss_cdas_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_wr_ss_cdas_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_maskcntl_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_ahb_defs_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/asib_ahbs/verilog/nic400_asib_ahbs_decode_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/amib_axim/verilog/nic400_amib_axim_undefs_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/amib_axim/verilog/nic400_amib_axim_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/amib_axim/verilog/nic400_amib_axim_chan_slice_hxb32.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/amib_axim/verilog/nic400_amib_axim_defs_hxb32.v"
`include "ips/nic400_hxb32/logical/nic400_hxb32/amib_axim/verilog/Ahb.v"
//`include "ips/nic400_hxb32/logical/nic400_hxb32/amib_axim/verilog/Ahb_undefs.v"
`include "modules/amba/rtl/ahb_axi_bdg.sv"
