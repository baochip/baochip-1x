// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

`include "modules/common/rtl/io_interface_def.sv"
`include "modules/common/rtl/amba_interface_def.sv"
`include "modules/common/rtl/ahbsramc.sv"
`include "modules/ifsub/rtl/ifsub1_intf.sv"
`include "modules/ifsub/rtl/udma_sub.sv"
`include "ips/L2_tcdm_hybrid_interco/RTL/lint_2_axi.sv"
`include "ips/udma/udma_camera/rtl/generic_mult8x8.sv"
`include "ips/udma/udma_camera/rtl/camera_if.sv"
`include "ips/udma/udma_camera/rtl/camera_reg_if.sv"
`include "ips/udma/udma_core/rtl/common/io_tx_fifo_dc.sv"
`include "ips/udma/udma_core/rtl/common/io_shiftreg.sv"
`include "ips/udma/udma_core/rtl/common/io_tx_fifo_mark.sv"
`include "ips/udma/udma_core/rtl/common/udma_ctrl.sv"
`include "ips/udma/udma_core/rtl/common/io_generic_fifo.sv"
`include "ips/udma/udma_core/rtl/common/io_event_counter.sv"
`include "ips/udma/udma_core/rtl/common/udma_clk_div_cnt.sv"
`include "ips/udma/udma_core/rtl/common/udma_apb4k_if.sv"
`include "ips/udma/udma_core/rtl/common/udma_dc_fifo.sv"
//`include "ips/udma/udma_core/rtl/common/io_clk_gen.sv"
`include "ips/udma/udma_core/rtl/common/io_tx_fifo.sv"
`include "ips/udma/udma_core/rtl/common/udma_clkgen.sv"
`include "ips/udma/udma_core/rtl/core/udma_rx_channels.sv"
`include "ips/udma/udma_core/rtl/core/udma_tx_channels.sv"
`include "ips/udma/udma_core/rtl/core/udma_core4k.sv"
`include "ips/udma/udma_core/rtl/core/udma_arbiter.sv"
`include "ips/udma/udma_core/rtl/core/udma_ch_addrgen.sv"
`include "ips/udma/udma_core/rtl/core/udma_stream_unit.sv"
`include "ips/udma/udma_external_per/rtl/udma_external_per_wrapper.sv"
`include "ips/udma/udma_external_per/rtl/udma_external_per_reg_if.sv"
`include "ips/udma/udma_external_per/rtl/udma_external_per_top.sv"
`include "ips/udma/udma_external_per/rtl/udma_traffic_gen_tx.sv"
`include "ips/udma/udma_external_per/rtl/udma_traffic_gen_rx.sv"
`include "ips/udma/udma_filter/rtl/udma_filter_au.sv"
`include "ips/udma/udma_filter/rtl/udma_filter_rx_dataout.sv"
`include "ips/udma/udma_filter/rtl/udma_filter_tx_datafetch.sv"
`include "ips/udma/udma_filter/rtl/udma_filter_reg_if.sv"
`include "ips/udma/udma_filter/rtl/udma_filter.sv"
`include "ips/udma/udma_filter/rtl/udma_filter_bincu.sv"
//`include "ips/udma/udma_i2c/rtl/udma_i2c_reg_if.sv"
//`include "ips/udma/udma_i2c/rtl/udma_i2c_bus_ctrl.sv"
//`include "ips/udma/udma_i2c/rtl/udma_i2c_top.sv"
//`include "ips/udma/udma_i2c/rtl/udma_i2c_control.sv"

`include "ips/udma/udma_i2c/rtl/udma_i2c_bus_ctrl.sv"
`include "ips/udma/udma_i2c/rtl/udma_i2c_control.sv"
`include "ips/udma/udma_i2c/rtl/udma_i2c_reg_if.sv"
`include "ips/udma/udma_i2c/rtl/udma_i2c_top.sv"
`include "ips/udma/udma_i2c/rtl/udma_i2c_undef.sv"


`include "ips/udma/udma_i2s/rtl/udma_i2s_top.sv"
`include "ips/udma/udma_i2s/rtl/i2s_txrx.sv"
`include "ips/udma/udma_i2s/rtl/i2s_clk_gen.sv"
`include "ips/udma/udma_i2s/rtl/i2s_clkws_gen.sv"
`include "ips/udma/udma_i2s/rtl/cic_top.sv"
`include "ips/udma/udma_i2s/rtl/i2s_tx_channel.sv"
`include "ips/udma/udma_i2s/rtl/pdm_top.sv"
`include "ips/udma/udma_i2s/rtl/udma_i2s_reg_if.sv"
`include "ips/udma/udma_i2s/rtl/i2s_rx_channel.sv"
`include "ips/udma/udma_i2s/rtl/cic_integrator.sv"
`include "ips/udma/udma_i2s/rtl/cic_comb.sv"
`include "ips/udma/udma_i2s/rtl/i2s_ws_gen.sv"
`include "ips/udma/udma_qspi/rtl/udma_spim_reg_if.sv"
`include "ips/udma/udma_qspi/rtl/udma_spim_top.sv"
`include "ips/udma/udma_qspi/rtl/udma_spim_ctrl.sv"
`include "ips/udma/udma_qspi/rtl/udma_spim_txrx.sv"
`include "ips/udma/udma_qspi/rtl/udma_spim_undef.sv"
`include "ips/udma/udma_sdio/rtl/sdio_txrx.sv"
`include "ips/udma/udma_sdio/rtl/sdio_crc7.sv"
`include "ips/udma/udma_sdio/rtl/udma_sdio_top.sv"
`include "ips/udma/udma_sdio/rtl/udma_sdio_reg_if.sv"
`include "ips/udma/udma_sdio/rtl/sdio_crc16.sv"
`include "ips/udma/udma_sdio/rtl/sdio_txrx_cmd.sv"
`include "ips/udma/udma_sdio/rtl/sdio_txrx_data.sv"
`include "ips/udma/udma_uart/rtl/udma_uart_tx.sv"
`include "ips/udma/udma_uart/rtl/udma_uart_reg_if.sv"
`include "ips/udma/udma_uart/rtl/udma_uart_rx.sv"
`include "ips/udma/udma_uart/rtl/udma_uart_top.sv"
`include "ips/axi/axi_slice_dc/src/dc_token_ring_fifo_din.v"
`include "ips/axi/axi_slice_dc/src/dc_token_ring_fifo_dout.v"
`include "ips/common_cells/src/deprecated/pulp_sync_wedge.sv"
`include "ips/tech_cells_generic/src/deprecated/pulp_clock_gating_async.sv"
`include "ips/tech_cells_generic/src/deprecated/pulp_clk_cells.sv"
`include "ips/axi/axi_slice_dc/src/dc_data_buffer.sv"
`include "ips/axi/axi_slice_dc/src/dc_full_detector.v"
`include "ips/axi/axi_slice_dc/src/dc_token_ring.v"
`include "ips/axi/axi_slice_dc/src/dc_synchronizer.v"
`include "ips/common_cells/src/deprecated/pulp_sync.sv"
`include "ips/common_cells/src/edge_propagator_rx.sv"
`include "ips/common_cells/src/edge_propagator.sv"
`include "ips/common_cells/src/edge_propagator_tx.sv"
`include "ips/common_cells/src/edge_propagator_ack.sv"
`include "ips/common_cells/src/onehot_to_bin.sv"
`include "modules/ifsub/rtl/udma_scif_reg.sv"
`include "modules/ifsub/rtl/udma_scif_rx.sv"
`include "modules/ifsub/rtl/udma_scif_tx.sv"
`include "modules/ifsub/rtl/udma_scif.sv"
`include "modules/ifsub/rtl/udma_spis_txrx.sv"
`include "modules/ifsub/rtl/udma_spis_reg.sv"
`include "modules/ifsub/rtl/udma_spis.sv"
//`include "rtl/common/icg_v0.2.v"
`include "modules/ifsub/rtl/iox.sv"
`include "modules/ifsub/rtl/pwm_intf.sv"
`include "modules/ifsub/rtl/udma_adc_ts_top.sv"
`include "modules/ifsub/rtl/udma_adc_ts_reg_if.sv"
`include "ips/apb/apb_adv_timer/rtl/adv_timer_apb_if.sv"
`include "ips/apb/apb_adv_timer/rtl/apb_adv_timer.sv"
`include "ips/apb/apb_adv_timer/rtl/comparator.sv"
`include "ips/apb/apb_adv_timer/rtl/input_stage.sv"
`include "ips/apb/apb_adv_timer/rtl/lut_4x4.sv"
`include "ips/apb/apb_adv_timer/rtl/out_filter.sv"
`include "ips/apb/apb_adv_timer/rtl/prescaler.sv"
`include "ips/apb/apb_adv_timer/rtl/timer_cntrl.sv"
`include "ips/apb/apb_adv_timer/rtl/timer_module.sv"
`include "ips/apb/apb_adv_timer/rtl/up_down_counter.sv"

`include "ips/ahb_bmxif2/ahb_bmxif_default_slave.v"
`include "ips/ahb_bmxif2/ahb_bmxif_intf.sv"
`include "ips/ahb_bmxif2/ahb_bmxif_lite.v"
`include "ips/ahb_bmxif2/ahb_bmxif.v"
`include "ips/ahb_bmxif2/ifabm0.v"
`include "ips/ahb_bmxif2/ifabm1.v"
`include "ips/ahb_bmxif2/ifabm2.v"
`include "ips/ahb_bmxif2/ifib.v"
`include "ips/ahb_bmxif2/ifmbs0.v"
`include "ips/ahb_bmxif2/ifmbs1.v"
`include "ips/ahb_bmxif2/ifmbs2.v"
`include "ips/ahb_bmxif2/ifobm0.v"
`include "ips/ahb_bmxif2/ifobm1.v"
`include "ips/ahb_bmxif2/ifobm2.v"
`ifdef SIM
`define ARM_UD_MODEL
`define ARM_DISABLE_EMA_CHECK
`include "asic_top/lib/arm_sram_macro/ifram32kx36/ifram32kx36.v"
`endif
`include "modules/ifsub/rtl/ifram.sv"

`include "modules/ifsub/rtl/soc_ifsub.sv"
`include "include/udc_inc.sv"
//`include "rtl/include/sddc_inc_v0.1.sv"
`include "include/bio_inc.sv"
