// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

`include "modules/dft/rtl/bscell.sv"
//`include "rtl/dft/jtag_enable.sv"
//`include "rtl/dft/jtag_enable_synch.sv"
`include "modules/dft/rtl/jtagreg.sv"
//`include "rtl/dft/jtag_rst_synch.sv"
`include "modules/dft/rtl/jtag_sync.sv"
`include "modules/dft/rtl/tap_top.sv"
`include "modules/dft/rtl/jtagtap.sv"