// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

`include "ips/pl230_udma/verilog/pl230_ahb_ctrl.v"
`include "ips/pl230_udma/verilog/pl230_apb_regs.v"
`include "ips/pl230_udma/verilog/pl230_dma_data.v"
`include "ips/pl230_udma/verilog/pl230_udma.v"

`include "modules/core/rtl/mdma.sv"