// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

//  Description : Toplevel Testbench Package
//                including all supporting modules/packages/tasks/functions
//
/////////////////////////////////////////////////////////////////////////// 


`include "tb_util_pkg.sv"
`include "daric_defs.sv"
`include "axi_tb_pkg.sv"
`include "axi_util_pkg.sv"
`include "ahb_tb_pkg.sv"
`include "ahb_tb_mst.sv"
`include "ahb_tb_mon.sv"
`include "axi_if_mst.sv"
`include "axi_if_bfm.sv"
`include "W25Q128JVxIM.v"
`include "W959D8NFYA.vcs.vp"
`include "i2cSlaveModules.v"
`include "iis_emu.sv"
`include "sdio_emu.sv"
`include "camera_emu.sv"
`include "usb_phy.sv"
`include "usb_host_emu.sv"
