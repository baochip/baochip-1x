// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

// Post-processing pass by bist_insert.py on 2025-02-08 04:21:34.811410

// -----------------------------------------------------------------------------
// Auto-Generated by:        __   _ __      _  __
//                          / /  (_) /____ | |/_/
//                         / /__/ / __/ -_)>  <
//                        /____/_/\__/\__/_/|_|
//                     Build your hardware, easily!
//                   https://github.com/enjoy-digital/litex
//
// Filename   : cram_axi.v
// Device     : 
// LiteX sha1 : 5375731c
// Date       : 2025-02-08 04:21:32
//------------------------------------------------------------------------------

`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// Module
//------------------------------------------------------------------------------

module cram_axi (
	rbif.slavedp	rbif_rdram1kx32[0:5],
	rbif.slavedp	rbif_rdram128x22[0:7],
	rbif.slavedp	rbif_rdram512x64[0:3],
    input  wire          aclk,
    input  wire          rst,
    input  wire          always_on,
    input  wire   [31:0] trimming_reset,
    input  wire          trimming_reset_ena,
    output wire          ibus_axi_awvalid,
    input  wire          ibus_axi_awready,
    output wire   [31:0] ibus_axi_awaddr,
    output wire    [1:0] ibus_axi_awburst,
    output wire    [7:0] ibus_axi_awlen,
    output wire    [2:0] ibus_axi_awsize,
    output wire          ibus_axi_awlock,
    output wire    [2:0] ibus_axi_awprot,
    output wire    [3:0] ibus_axi_awcache,
    output wire    [3:0] ibus_axi_awqos,
    output wire    [3:0] ibus_axi_awregion,
    output wire          ibus_axi_awid,
    output wire          ibus_axi_awuser,
    output wire          ibus_axi_wvalid,
    input  wire          ibus_axi_wready,
    output wire          ibus_axi_wlast,
    output wire   [63:0] ibus_axi_wdata,
    output wire    [7:0] ibus_axi_wstrb,
    output wire          ibus_axi_wuser,
    input  wire          ibus_axi_bvalid,
    output wire          ibus_axi_bready,
    input  wire    [1:0] ibus_axi_bresp,
    input  wire          ibus_axi_bid,
    input  wire          ibus_axi_buser,
    output wire          ibus_axi_arvalid,
    input  wire          ibus_axi_arready,
    output wire   [31:0] ibus_axi_araddr,
    output wire    [1:0] ibus_axi_arburst,
    output wire    [7:0] ibus_axi_arlen,
    output wire    [2:0] ibus_axi_arsize,
    output wire          ibus_axi_arlock,
    output wire    [2:0] ibus_axi_arprot,
    output wire    [3:0] ibus_axi_arcache,
    output wire    [3:0] ibus_axi_arqos,
    output wire    [3:0] ibus_axi_arregion,
    output wire          ibus_axi_arid,
    output wire          ibus_axi_aruser,
    input  wire          ibus_axi_rvalid,
    output wire          ibus_axi_rready,
    input  wire          ibus_axi_rlast,
    input  wire    [1:0] ibus_axi_rresp,
    input  wire   [63:0] ibus_axi_rdata,
    input  wire          ibus_axi_rid,
    input  wire          ibus_axi_ruser,
    output wire          dbus_axi_awvalid,
    input  wire          dbus_axi_awready,
    output wire   [31:0] dbus_axi_awaddr,
    output wire    [1:0] dbus_axi_awburst,
    output wire    [7:0] dbus_axi_awlen,
    output wire    [2:0] dbus_axi_awsize,
    output wire          dbus_axi_awlock,
    output wire    [2:0] dbus_axi_awprot,
    output wire    [3:0] dbus_axi_awcache,
    output wire    [3:0] dbus_axi_awqos,
    output wire    [3:0] dbus_axi_awregion,
    output wire          dbus_axi_awid,
    output wire          dbus_axi_awuser,
    output wire          dbus_axi_wvalid,
    input  wire          dbus_axi_wready,
    output wire          dbus_axi_wlast,
    output wire   [31:0] dbus_axi_wdata,
    output wire    [3:0] dbus_axi_wstrb,
    output wire          dbus_axi_wuser,
    input  wire          dbus_axi_bvalid,
    output wire          dbus_axi_bready,
    input  wire    [1:0] dbus_axi_bresp,
    input  wire          dbus_axi_bid,
    input  wire          dbus_axi_buser,
    output wire          dbus_axi_arvalid,
    input  wire          dbus_axi_arready,
    output wire   [31:0] dbus_axi_araddr,
    output wire    [1:0] dbus_axi_arburst,
    output wire    [7:0] dbus_axi_arlen,
    output wire    [2:0] dbus_axi_arsize,
    output wire          dbus_axi_arlock,
    output wire    [2:0] dbus_axi_arprot,
    output wire    [3:0] dbus_axi_arcache,
    output wire    [3:0] dbus_axi_arqos,
    output wire    [3:0] dbus_axi_arregion,
    output wire          dbus_axi_arid,
    output wire          dbus_axi_aruser,
    input  wire          dbus_axi_rvalid,
    output wire          dbus_axi_rready,
    input  wire          dbus_axi_rlast,
    input  wire    [1:0] dbus_axi_rresp,
    input  wire   [31:0] dbus_axi_rdata,
    input  wire          dbus_axi_rid,
    input  wire          dbus_axi_ruser,
    output wire          p_axi_awvalid,
    input  wire          p_axi_awready,
    output wire   [31:0] p_axi_awaddr,
    output wire    [2:0] p_axi_awprot,
    output wire          p_axi_wvalid,
    input  wire          p_axi_wready,
    output wire   [31:0] p_axi_wdata,
    output wire    [3:0] p_axi_wstrb,
    input  wire          p_axi_bvalid,
    output wire          p_axi_bready,
    input  wire    [1:0] p_axi_bresp,
    output wire          p_axi_arvalid,
    input  wire          p_axi_arready,
    output wire   [31:0] p_axi_araddr,
    output wire    [2:0] p_axi_arprot,
    input  wire          p_axi_rvalid,
    output wire          p_axi_rready,
    input  wire    [1:0] p_axi_rresp,
    input  wire   [31:0] p_axi_rdata,
    input  wire          jtag_tdi,
    output wire          jtag_tdo,
    input  wire          jtag_tms,
    input  wire          jtag_tck,
    input  wire          jtag_trst_n,
    input  wire          cmbist,
    input  wire          cmatpg,
    input  wire    [2:0] vexsramtrm,
    output reg     [7:0] coreuser_vex,
    output reg           vex_mm,
    input  wire    [1:0] default_user,
    input  wire          default_mm,
    output wire          sleep_req,
    input  wire   [15:0] irqarray_bank0,
    input  wire   [15:0] irqarray_bank1,
    input  wire   [15:0] irqarray_bank2,
    input  wire   [15:0] irqarray_bank3,
    input  wire   [15:0] irqarray_bank4,
    input  wire   [15:0] irqarray_bank5,
    input  wire   [15:0] irqarray_bank6,
    input  wire   [15:0] irqarray_bank7,
    input  wire   [15:0] irqarray_bank8,
    input  wire   [15:0] irqarray_bank9,
    input  wire   [15:0] irqarray_bank10,
    input  wire   [15:0] irqarray_bank11,
    input  wire   [15:0] irqarray_bank12,
    input  wire   [15:0] irqarray_bank13,
    input  wire   [15:0] irqarray_bank14,
    input  wire   [15:0] irqarray_bank15,
    input  wire   [15:0] irqarray_bank16,
    input  wire   [15:0] irqarray_bank17,
    input  wire   [15:0] irqarray_bank18,
    input  wire   [15:0] irqarray_bank19,
    input  wire   [31:0] mbox_w_dat,
    input  wire          mbox_w_valid,
    output wire          mbox_w_ready,
    input  wire          mbox_w_done,
    output wire   [31:0] mbox_r_dat,
    output wire          mbox_r_valid,
    input  wire          mbox_r_ready,
    output wire          mbox_r_done,
    input  wire          mbox_w_abort,
    output wire          mbox_r_abort,
    output wire   [31:0] test
);


//------------------------------------------------------------------------------
// Signals
//------------------------------------------------------------------------------

wire          sys_clk;
wire          sys_rst;
wire          always_on_clk;
wire          always_on_rst;
reg    [31:0] cramsoc_interrupt;
wire   [31:0] cramsoc_trimming_reset;
wire          cramsoc_trimming_reset_ena;
wire          cramsoc_satp_mode;
wire    [8:0] cramsoc_satp_asid;
wire   [21:0] cramsoc_satp_ppn;
wire          cramsoc_wfi_active;
wire    [1:0] cramsoc_privilege;
wire          cramsoc_cmbist;
wire          cramsoc_cmatpg;
wire    [2:0] cramsoc_vexsramtrm;
reg           cramsoc_ibus_axi_aw_valid;
wire          cramsoc_ibus_axi_aw_ready;
reg    [31:0] cramsoc_ibus_axi_aw_payload_addr;
reg     [1:0] cramsoc_ibus_axi_aw_payload_burst;
reg     [7:0] cramsoc_ibus_axi_aw_payload_len;
reg     [2:0] cramsoc_ibus_axi_aw_payload_size;
reg           cramsoc_ibus_axi_aw_payload_lock;
reg     [2:0] cramsoc_ibus_axi_aw_payload_prot;
reg     [3:0] cramsoc_ibus_axi_aw_payload_cache;
reg     [3:0] cramsoc_ibus_axi_aw_payload_qos;
reg     [3:0] cramsoc_ibus_axi_aw_payload_region;
reg           cramsoc_ibus_axi_aw_param_id;
reg           cramsoc_ibus_axi_aw_param_user;
reg           cramsoc_ibus_axi_w_valid;
wire          cramsoc_ibus_axi_w_ready;
reg           cramsoc_ibus_axi_w_last;
reg    [63:0] cramsoc_ibus_axi_w_payload_data;
reg     [7:0] cramsoc_ibus_axi_w_payload_strb;
reg           cramsoc_ibus_axi_w_param_user;
wire          cramsoc_ibus_axi_b_valid;
reg           cramsoc_ibus_axi_b_ready;
wire    [1:0] cramsoc_ibus_axi_b_payload_resp;
wire          cramsoc_ibus_axi_b_param_id;
wire          cramsoc_ibus_axi_b_param_user;
wire          cramsoc_ibus_axi_ar_valid;
wire          cramsoc_ibus_axi_ar_ready;
wire   [31:0] cramsoc_ibus_axi_ar_payload_addr;
wire    [1:0] cramsoc_ibus_axi_ar_payload_burst;
wire    [7:0] cramsoc_ibus_axi_ar_payload_len;
wire    [2:0] cramsoc_ibus_axi_ar_payload_size;
wire          cramsoc_ibus_axi_ar_payload_lock;
wire    [2:0] cramsoc_ibus_axi_ar_payload_prot;
wire    [3:0] cramsoc_ibus_axi_ar_payload_cache;
wire    [3:0] cramsoc_ibus_axi_ar_payload_qos;
wire    [3:0] cramsoc_ibus_axi_ar_payload_region;
wire          cramsoc_ibus_axi_ar_param_id;
reg           cramsoc_ibus_axi_ar_param_user;
wire          cramsoc_ibus_axi_r_valid;
wire          cramsoc_ibus_axi_r_ready;
wire          cramsoc_ibus_axi_r_last;
wire    [1:0] cramsoc_ibus_axi_r_payload_resp;
wire   [63:0] cramsoc_ibus_axi_r_payload_data;
wire          cramsoc_ibus_axi_r_param_id;
wire          cramsoc_ibus_axi_r_param_user;
wire          cramsoc_dbus_axi_aw_valid;
wire          cramsoc_dbus_axi_aw_ready;
wire   [31:0] cramsoc_dbus_axi_aw_payload_addr;
wire    [1:0] cramsoc_dbus_axi_aw_payload_burst;
wire    [7:0] cramsoc_dbus_axi_aw_payload_len;
wire    [2:0] cramsoc_dbus_axi_aw_payload_size;
wire          cramsoc_dbus_axi_aw_payload_lock;
wire    [2:0] cramsoc_dbus_axi_aw_payload_prot;
wire    [3:0] cramsoc_dbus_axi_aw_payload_cache;
wire    [3:0] cramsoc_dbus_axi_aw_payload_qos;
wire    [3:0] cramsoc_dbus_axi_aw_payload_region;
wire          cramsoc_dbus_axi_aw_param_id;
reg           cramsoc_dbus_axi_aw_param_user;
wire          cramsoc_dbus_axi_w_valid;
wire          cramsoc_dbus_axi_w_ready;
wire          cramsoc_dbus_axi_w_last;
wire   [31:0] cramsoc_dbus_axi_w_payload_data;
wire    [3:0] cramsoc_dbus_axi_w_payload_strb;
reg           cramsoc_dbus_axi_w_param_user;
wire          cramsoc_dbus_axi_b_valid;
wire          cramsoc_dbus_axi_b_ready;
wire    [1:0] cramsoc_dbus_axi_b_payload_resp;
wire          cramsoc_dbus_axi_b_param_id;
wire          cramsoc_dbus_axi_b_param_user;
wire          cramsoc_dbus_axi_ar_valid;
wire          cramsoc_dbus_axi_ar_ready;
wire   [31:0] cramsoc_dbus_axi_ar_payload_addr;
wire    [1:0] cramsoc_dbus_axi_ar_payload_burst;
wire    [7:0] cramsoc_dbus_axi_ar_payload_len;
wire    [2:0] cramsoc_dbus_axi_ar_payload_size;
wire          cramsoc_dbus_axi_ar_payload_lock;
wire    [2:0] cramsoc_dbus_axi_ar_payload_prot;
wire    [3:0] cramsoc_dbus_axi_ar_payload_cache;
wire    [3:0] cramsoc_dbus_axi_ar_payload_qos;
wire    [3:0] cramsoc_dbus_axi_ar_payload_region;
wire          cramsoc_dbus_axi_ar_param_id;
reg           cramsoc_dbus_axi_ar_param_user;
wire          cramsoc_dbus_axi_r_valid;
wire          cramsoc_dbus_axi_r_ready;
wire          cramsoc_dbus_axi_r_last;
wire    [1:0] cramsoc_dbus_axi_r_payload_resp;
wire   [31:0] cramsoc_dbus_axi_r_payload_data;
wire          cramsoc_dbus_axi_r_param_id;
wire          cramsoc_dbus_axi_r_param_user;
wire          cramsoc_dbus_peri_aw_valid;
wire          cramsoc_dbus_peri_aw_ready;
wire   [31:0] cramsoc_dbus_peri_aw_payload_addr;
wire    [1:0] cramsoc_dbus_peri_aw_payload_burst;
wire    [7:0] cramsoc_dbus_peri_aw_payload_len;
wire    [2:0] cramsoc_dbus_peri_aw_payload_size;
wire          cramsoc_dbus_peri_aw_payload_lock;
wire    [2:0] cramsoc_dbus_peri_aw_payload_prot;
wire    [3:0] cramsoc_dbus_peri_aw_payload_cache;
wire    [3:0] cramsoc_dbus_peri_aw_payload_qos;
wire    [3:0] cramsoc_dbus_peri_aw_payload_region;
wire          cramsoc_dbus_peri_aw_param_id;
wire          cramsoc_dbus_peri_aw_param_user;
wire          cramsoc_dbus_peri_w_valid;
wire          cramsoc_dbus_peri_w_ready;
wire          cramsoc_dbus_peri_w_last;
wire   [31:0] cramsoc_dbus_peri_w_payload_data;
wire    [3:0] cramsoc_dbus_peri_w_payload_strb;
wire          cramsoc_dbus_peri_w_param_user;
wire          cramsoc_dbus_peri_b_valid;
wire          cramsoc_dbus_peri_b_ready;
wire    [1:0] cramsoc_dbus_peri_b_payload_resp;
wire          cramsoc_dbus_peri_b_param_id;
reg           cramsoc_dbus_peri_b_param_user;
wire          cramsoc_dbus_peri_ar_valid;
wire          cramsoc_dbus_peri_ar_ready;
wire   [31:0] cramsoc_dbus_peri_ar_payload_addr;
wire    [1:0] cramsoc_dbus_peri_ar_payload_burst;
wire    [7:0] cramsoc_dbus_peri_ar_payload_len;
wire    [2:0] cramsoc_dbus_peri_ar_payload_size;
wire          cramsoc_dbus_peri_ar_payload_lock;
wire    [2:0] cramsoc_dbus_peri_ar_payload_prot;
wire    [3:0] cramsoc_dbus_peri_ar_payload_cache;
wire    [3:0] cramsoc_dbus_peri_ar_payload_qos;
wire    [3:0] cramsoc_dbus_peri_ar_payload_region;
wire          cramsoc_dbus_peri_ar_param_id;
wire          cramsoc_dbus_peri_ar_param_user;
wire          cramsoc_dbus_peri_r_valid;
wire          cramsoc_dbus_peri_r_ready;
wire          cramsoc_dbus_peri_r_last;
wire    [1:0] cramsoc_dbus_peri_r_payload_resp;
wire   [31:0] cramsoc_dbus_peri_r_payload_data;
wire          cramsoc_dbus_peri_r_param_id;
reg           cramsoc_dbus_peri_r_param_user;
wire          cramsoc_peripherals_aw_valid;
wire          cramsoc_peripherals_aw_ready;
wire   [31:0] cramsoc_peripherals_aw_payload_addr;
wire    [2:0] cramsoc_peripherals_aw_payload_prot;
wire          cramsoc_peripherals_w_valid;
wire          cramsoc_peripherals_w_ready;
wire   [31:0] cramsoc_peripherals_w_payload_data;
wire    [3:0] cramsoc_peripherals_w_payload_strb;
wire          cramsoc_peripherals_b_valid;
wire          cramsoc_peripherals_b_ready;
wire    [1:0] cramsoc_peripherals_b_payload_resp;
wire          cramsoc_peripherals_ar_valid;
wire          cramsoc_peripherals_ar_ready;
wire   [31:0] cramsoc_peripherals_ar_payload_addr;
wire    [2:0] cramsoc_peripherals_ar_payload_prot;
wire          cramsoc_peripherals_r_valid;
wire          cramsoc_peripherals_r_ready;
wire    [1:0] cramsoc_peripherals_r_payload_resp;
wire   [31:0] cramsoc_peripherals_r_payload_data;
wire          cramsoc_axi_csr_aw_valid;
wire          cramsoc_axi_csr_aw_ready;
wire   [31:0] cramsoc_axi_csr_aw_payload_addr;
wire    [1:0] cramsoc_axi_csr_aw_payload_burst;
wire    [7:0] cramsoc_axi_csr_aw_payload_len;
wire    [2:0] cramsoc_axi_csr_aw_payload_size;
wire          cramsoc_axi_csr_aw_payload_lock;
wire    [2:0] cramsoc_axi_csr_aw_payload_prot;
wire    [3:0] cramsoc_axi_csr_aw_payload_cache;
wire    [3:0] cramsoc_axi_csr_aw_payload_qos;
wire    [3:0] cramsoc_axi_csr_aw_payload_region;
wire          cramsoc_axi_csr_aw_param_id;
wire          cramsoc_axi_csr_aw_param_user;
wire          cramsoc_axi_csr_w_valid;
wire          cramsoc_axi_csr_w_ready;
wire          cramsoc_axi_csr_w_last;
wire   [31:0] cramsoc_axi_csr_w_payload_data;
wire    [3:0] cramsoc_axi_csr_w_payload_strb;
wire          cramsoc_axi_csr_w_param_user;
wire          cramsoc_axi_csr_b_valid;
wire          cramsoc_axi_csr_b_ready;
wire    [1:0] cramsoc_axi_csr_b_payload_resp;
wire          cramsoc_axi_csr_b_param_id;
reg           cramsoc_axi_csr_b_param_user;
wire          cramsoc_axi_csr_ar_valid;
wire          cramsoc_axi_csr_ar_ready;
wire   [31:0] cramsoc_axi_csr_ar_payload_addr;
wire    [1:0] cramsoc_axi_csr_ar_payload_burst;
wire    [7:0] cramsoc_axi_csr_ar_payload_len;
wire    [2:0] cramsoc_axi_csr_ar_payload_size;
wire          cramsoc_axi_csr_ar_payload_lock;
wire    [2:0] cramsoc_axi_csr_ar_payload_prot;
wire    [3:0] cramsoc_axi_csr_ar_payload_cache;
wire    [3:0] cramsoc_axi_csr_ar_payload_qos;
wire    [3:0] cramsoc_axi_csr_ar_payload_region;
wire          cramsoc_axi_csr_ar_param_id;
wire          cramsoc_axi_csr_ar_param_user;
wire          cramsoc_axi_csr_r_valid;
wire          cramsoc_axi_csr_r_ready;
wire          cramsoc_axi_csr_r_last;
wire    [1:0] cramsoc_axi_csr_r_payload_resp;
wire   [31:0] cramsoc_axi_csr_r_payload_data;
wire          cramsoc_axi_csr_r_param_id;
reg           cramsoc_axi_csr_r_param_user;
wire          cramsoc_corecsr_aw_valid;
wire          cramsoc_corecsr_aw_ready;
reg           cramsoc_corecsr_aw_first;
reg           cramsoc_corecsr_aw_last;
wire   [31:0] cramsoc_corecsr_aw_payload_addr;
wire    [2:0] cramsoc_corecsr_aw_payload_prot;
wire          cramsoc_corecsr_w_valid;
wire          cramsoc_corecsr_w_ready;
reg           cramsoc_corecsr_w_first;
reg           cramsoc_corecsr_w_last;
wire   [31:0] cramsoc_corecsr_w_payload_data;
wire    [3:0] cramsoc_corecsr_w_payload_strb;
wire          cramsoc_corecsr_b_valid;
wire          cramsoc_corecsr_b_ready;
wire          cramsoc_corecsr_b_first;
wire          cramsoc_corecsr_b_last;
wire    [1:0] cramsoc_corecsr_b_payload_resp;
wire          cramsoc_corecsr_ar_valid;
wire          cramsoc_corecsr_ar_ready;
reg           cramsoc_corecsr_ar_first;
reg           cramsoc_corecsr_ar_last;
wire   [31:0] cramsoc_corecsr_ar_payload_addr;
wire    [2:0] cramsoc_corecsr_ar_payload_prot;
wire          cramsoc_corecsr_r_valid;
wire          cramsoc_corecsr_r_ready;
wire          cramsoc_corecsr_r_first;
wire          cramsoc_corecsr_r_last;
wire    [1:0] cramsoc_corecsr_r_payload_resp;
wire   [31:0] cramsoc_corecsr_r_payload_data;
wire          cramsoc_dbus_aw_valid;
wire          cramsoc_dbus_aw_ready;
wire   [31:0] cramsoc_dbus_aw_payload_addr;
wire    [1:0] cramsoc_dbus_aw_payload_burst;
wire    [7:0] cramsoc_dbus_aw_payload_len;
wire    [2:0] cramsoc_dbus_aw_payload_size;
wire          cramsoc_dbus_aw_payload_lock;
wire    [2:0] cramsoc_dbus_aw_payload_prot;
wire    [3:0] cramsoc_dbus_aw_payload_cache;
wire    [3:0] cramsoc_dbus_aw_payload_qos;
wire    [3:0] cramsoc_dbus_aw_payload_region;
wire          cramsoc_dbus_aw_param_id;
wire          cramsoc_dbus_aw_param_user;
wire          cramsoc_dbus_w_valid;
wire          cramsoc_dbus_w_ready;
wire          cramsoc_dbus_w_last;
wire   [31:0] cramsoc_dbus_w_payload_data;
wire    [3:0] cramsoc_dbus_w_payload_strb;
wire          cramsoc_dbus_w_param_user;
wire          cramsoc_dbus_b_valid;
wire          cramsoc_dbus_b_ready;
wire    [1:0] cramsoc_dbus_b_payload_resp;
wire          cramsoc_dbus_b_param_id;
wire          cramsoc_dbus_b_param_user;
wire          cramsoc_dbus_ar_valid;
wire          cramsoc_dbus_ar_ready;
wire   [31:0] cramsoc_dbus_ar_payload_addr;
wire    [1:0] cramsoc_dbus_ar_payload_burst;
wire    [7:0] cramsoc_dbus_ar_payload_len;
wire    [2:0] cramsoc_dbus_ar_payload_size;
wire          cramsoc_dbus_ar_payload_lock;
wire    [2:0] cramsoc_dbus_ar_payload_prot;
wire    [3:0] cramsoc_dbus_ar_payload_cache;
wire    [3:0] cramsoc_dbus_ar_payload_qos;
wire    [3:0] cramsoc_dbus_ar_payload_region;
wire          cramsoc_dbus_ar_param_id;
wire          cramsoc_dbus_ar_param_user;
wire          cramsoc_dbus_r_valid;
wire          cramsoc_dbus_r_ready;
wire          cramsoc_dbus_r_last;
wire    [1:0] cramsoc_dbus_r_payload_resp;
wire   [31:0] cramsoc_dbus_r_payload_data;
wire          cramsoc_dbus_r_param_id;
wire          cramsoc_dbus_r_param_user;
reg    [31:0] cramsoc_vexriscvaxi_reset_mux;
reg    [31:0] cramsoc_vexriscvaxi;
reg    [31:0] cramsoc_load_storage;
reg           cramsoc_load_re;
reg    [31:0] cramsoc_reload_storage;
reg           cramsoc_reload_re;
reg           cramsoc_en_storage;
reg           cramsoc_en_re;
reg           cramsoc_update_value_storage;
reg           cramsoc_update_value_re;
reg    [31:0] cramsoc_value_status;
wire          cramsoc_value_we;
reg           cramsoc_value_re;
wire          cramsoc_irq;
wire          cramsoc_zero_status;
reg           cramsoc_zero_pending;
wire          cramsoc_zero_trigger;
reg           cramsoc_zero_clear;
reg           cramsoc_zero_trigger_d;
wire          cramsoc_zero0;
wire          cramsoc_status_status;
wire          cramsoc_status_we;
reg           cramsoc_status_re;
wire          cramsoc_zero1;
wire          cramsoc_pending_status;
wire          cramsoc_pending_we;
reg           cramsoc_pending_re;
reg           cramsoc_pending_r;
wire          cramsoc_zero2;
reg           cramsoc_enable_storage;
reg           cramsoc_enable_re;
reg    [31:0] cramsoc_value;
wire          o_resetOut;
reg           reset_debug_logic;
reg           debug_reset;
wire   [31:0] trimming_reset_1;
wire          trimming_reset_ena_1;
wire   [31:0] status;
wire          we;
reg           re;
reg    [31:0] latched_value;
wire          coreuser_enable0;
wire          coreuser_invert_priv0;
reg     [1:0] coreuser_control_storage;
reg           coreuser_control_re;
reg     [7:0] coreuser_coreuser;
reg           coreuser_mm;
reg     [8:0] coreuser_status_status;
wire          coreuser_status_we;
reg           coreuser_status_re;
wire    [7:0] coreuser_lut00;
wire    [7:0] coreuser_lut10;
wire    [7:0] coreuser_lut20;
wire    [7:0] coreuser_lut30;
reg    [31:0] coreuser_map_lo_storage;
reg           coreuser_map_lo_re;
wire    [7:0] coreuser_lut40;
wire    [7:0] coreuser_lut50;
wire    [7:0] coreuser_lut60;
wire    [7:0] coreuser_lut70;
reg    [31:0] coreuser_map_hi_storage;
reg           coreuser_map_hi_re;
wire    [1:0] coreuser_user00;
wire    [1:0] coreuser_user10;
wire    [1:0] coreuser_user20;
wire    [1:0] coreuser_user30;
wire    [1:0] coreuser_user40;
wire    [1:0] coreuser_user50;
wire    [1:0] coreuser_user60;
wire    [1:0] coreuser_user70;
wire    [1:0] coreuser_default;
reg    [17:0] coreuser_uservalue_storage;
reg           coreuser_uservalue_re;
reg           coreuser_protect_storage;
reg           coreuser_protect_re;
wire          coreuser_protect;
reg           coreuser_enable1;
reg           coreuser_invert_priv1;
reg     [7:0] coreuser_lut01;
reg     [7:0] coreuser_lut11;
reg     [7:0] coreuser_lut21;
reg     [7:0] coreuser_lut31;
reg     [7:0] coreuser_lut41;
reg     [7:0] coreuser_lut51;
reg     [7:0] coreuser_lut61;
reg     [7:0] coreuser_lut71;
reg     [1:0] coreuser_user01;
reg     [1:0] coreuser_user11;
reg     [1:0] coreuser_user21;
reg     [1:0] coreuser_user31;
reg     [1:0] coreuser_user41;
reg     [1:0] coreuser_user51;
reg     [1:0] coreuser_user61;
reg     [1:0] coreuser_user71;
reg     [1:0] coreuser_user_default;
reg     [1:0] coreuser_coreuser_2bit;
reg     [3:0] coreuser_coreuser_4bit;
reg           cpu_int_active;
wire          axi_active;
reg           ibus_r_active;
reg           dbus_r_active;
reg           dbus_w_active;
reg           pbus_r_active;
reg           pbus_w_active;
reg     [6:0] active_timeout;
reg    [15:0] irq_remap0;
reg    [15:0] irq_remap1;
reg    [15:0] irq_remap2;
reg    [15:0] irq_remap3;
reg    [15:0] irq_remap4;
reg    [15:0] irq_remap5;
reg    [15:0] irq_remap6;
reg    [15:0] irq_remap7;
reg    [15:0] irq_remap8;
reg    [15:0] irq_remap9;
reg    [15:0] irq_remap10;
reg    [15:0] irq_remap11;
reg    [15:0] irq_remap12;
reg    [15:0] irq_remap13;
reg    [15:0] irq_remap14;
reg    [15:0] irq_remap15;
reg    [15:0] irq_remap16;
reg    [15:0] irq_remap17;
reg    [15:0] irq_remap18;
reg    [15:0] irq_remap19;
wire          irqarray0_irq;
wire   [15:0] irqarray0_interrupts;
reg    [15:0] irqarray0_trigger;
reg    [15:0] irqarray0_soft_storage;
reg           irqarray0_soft_re;
wire   [15:0] irqarray0_use_edge;
reg    [15:0] irqarray0_edge_triggered_storage;
reg           irqarray0_edge_triggered_re;
wire   [15:0] irqarray0_rising;
reg    [15:0] irqarray0_polarity_storage;
reg           irqarray0_polarity_re;
wire          irqarray0_eventsourceflex0_status;
reg           irqarray0_eventsourceflex0_pending;
reg           irqarray0_eventsourceflex0_clear;
reg           irqarray0_eventsourceflex0_trigger_d;
reg           irqarray0_eventsourceflex0_trigger_filtered;
wire          irqarray0_eventsourceflex1_status;
reg           irqarray0_eventsourceflex1_pending;
reg           irqarray0_eventsourceflex1_clear;
reg           irqarray0_eventsourceflex1_trigger_d;
reg           irqarray0_eventsourceflex1_trigger_filtered;
wire          irqarray0_eventsourceflex2_status;
reg           irqarray0_eventsourceflex2_pending;
reg           irqarray0_eventsourceflex2_clear;
reg           irqarray0_eventsourceflex2_trigger_d;
reg           irqarray0_eventsourceflex2_trigger_filtered;
wire          irqarray0_eventsourceflex3_status;
reg           irqarray0_eventsourceflex3_pending;
reg           irqarray0_eventsourceflex3_clear;
reg           irqarray0_eventsourceflex3_trigger_d;
reg           irqarray0_eventsourceflex3_trigger_filtered;
wire          irqarray0_eventsourceflex4_status;
reg           irqarray0_eventsourceflex4_pending;
reg           irqarray0_eventsourceflex4_clear;
reg           irqarray0_eventsourceflex4_trigger_d;
reg           irqarray0_eventsourceflex4_trigger_filtered;
wire          irqarray0_eventsourceflex5_status;
reg           irqarray0_eventsourceflex5_pending;
reg           irqarray0_eventsourceflex5_clear;
reg           irqarray0_eventsourceflex5_trigger_d;
reg           irqarray0_eventsourceflex5_trigger_filtered;
wire          irqarray0_eventsourceflex6_status;
reg           irqarray0_eventsourceflex6_pending;
reg           irqarray0_eventsourceflex6_clear;
reg           irqarray0_eventsourceflex6_trigger_d;
reg           irqarray0_eventsourceflex6_trigger_filtered;
wire          irqarray0_eventsourceflex7_status;
reg           irqarray0_eventsourceflex7_pending;
reg           irqarray0_eventsourceflex7_clear;
reg           irqarray0_eventsourceflex7_trigger_d;
reg           irqarray0_eventsourceflex7_trigger_filtered;
wire          irqarray0_eventsourceflex8_status;
reg           irqarray0_eventsourceflex8_pending;
reg           irqarray0_eventsourceflex8_clear;
reg           irqarray0_eventsourceflex8_trigger_d;
reg           irqarray0_eventsourceflex8_trigger_filtered;
wire          irqarray0_eventsourceflex9_status;
reg           irqarray0_eventsourceflex9_pending;
reg           irqarray0_eventsourceflex9_clear;
reg           irqarray0_eventsourceflex9_trigger_d;
reg           irqarray0_eventsourceflex9_trigger_filtered;
wire          irqarray0_eventsourceflex10_status;
reg           irqarray0_eventsourceflex10_pending;
reg           irqarray0_eventsourceflex10_clear;
reg           irqarray0_eventsourceflex10_trigger_d;
reg           irqarray0_eventsourceflex10_trigger_filtered;
wire          irqarray0_eventsourceflex11_status;
reg           irqarray0_eventsourceflex11_pending;
reg           irqarray0_eventsourceflex11_clear;
reg           irqarray0_eventsourceflex11_trigger_d;
reg           irqarray0_eventsourceflex11_trigger_filtered;
wire          irqarray0_eventsourceflex12_status;
reg           irqarray0_eventsourceflex12_pending;
reg           irqarray0_eventsourceflex12_clear;
reg           irqarray0_eventsourceflex12_trigger_d;
reg           irqarray0_eventsourceflex12_trigger_filtered;
wire          irqarray0_eventsourceflex13_status;
reg           irqarray0_eventsourceflex13_pending;
reg           irqarray0_eventsourceflex13_clear;
reg           irqarray0_eventsourceflex13_trigger_d;
reg           irqarray0_eventsourceflex13_trigger_filtered;
wire          irqarray0_eventsourceflex14_status;
reg           irqarray0_eventsourceflex14_pending;
reg           irqarray0_eventsourceflex14_clear;
reg           irqarray0_eventsourceflex14_trigger_d;
reg           irqarray0_eventsourceflex14_trigger_filtered;
wire          irqarray0_eventsourceflex15_status;
reg           irqarray0_eventsourceflex15_pending;
reg           irqarray0_eventsourceflex15_clear;
reg           irqarray0_eventsourceflex15_trigger_d;
reg           irqarray0_eventsourceflex15_trigger_filtered;
wire          irqarray0_mdmairq_dupe0;
wire          irqarray0_nc_b0s10;
wire          irqarray0_nc_b0s20;
wire          irqarray0_nc_b0s30;
wire          irqarray0_pioirq0_dupe0;
wire          irqarray0_pioirq1_dupe0;
wire          irqarray0_pioirq2_dupe0;
wire          irqarray0_pioirq3_dupe0;
wire          irqarray0_nc_b0s80;
wire          irqarray0_nc_b0s90;
wire          irqarray0_nc_b0s100;
wire          irqarray0_nc_b0s110;
wire          irqarray0_nc_b0s120;
wire          irqarray0_nc_b0s130;
wire          irqarray0_nc_b0s140;
wire          irqarray0_nc_b0s150;
reg    [15:0] irqarray0_status_status;
wire          irqarray0_status_we;
reg           irqarray0_status_re;
wire          irqarray0_mdmairq_dupe1;
wire          irqarray0_nc_b0s11;
wire          irqarray0_nc_b0s21;
wire          irqarray0_nc_b0s31;
wire          irqarray0_pioirq0_dupe1;
wire          irqarray0_pioirq1_dupe1;
wire          irqarray0_pioirq2_dupe1;
wire          irqarray0_pioirq3_dupe1;
wire          irqarray0_nc_b0s81;
wire          irqarray0_nc_b0s91;
wire          irqarray0_nc_b0s101;
wire          irqarray0_nc_b0s111;
wire          irqarray0_nc_b0s121;
wire          irqarray0_nc_b0s131;
wire          irqarray0_nc_b0s141;
wire          irqarray0_nc_b0s151;
reg    [15:0] irqarray0_pending_status;
wire          irqarray0_pending_we;
reg           irqarray0_pending_re;
reg    [15:0] irqarray0_pending_r;
wire          irqarray0_mdmairq_dupe2;
wire          irqarray0_nc_b0s12;
wire          irqarray0_nc_b0s22;
wire          irqarray0_nc_b0s32;
wire          irqarray0_pioirq0_dupe2;
wire          irqarray0_pioirq1_dupe2;
wire          irqarray0_pioirq2_dupe2;
wire          irqarray0_pioirq3_dupe2;
wire          irqarray0_nc_b0s82;
wire          irqarray0_nc_b0s92;
wire          irqarray0_nc_b0s102;
wire          irqarray0_nc_b0s112;
wire          irqarray0_nc_b0s122;
wire          irqarray0_nc_b0s132;
wire          irqarray0_nc_b0s142;
wire          irqarray0_nc_b0s152;
reg    [15:0] irqarray0_enable_storage;
reg           irqarray0_enable_re;
wire          irqarray1_irq;
wire   [15:0] irqarray1_interrupts;
reg    [15:0] irqarray1_trigger;
reg    [15:0] irqarray1_soft_storage;
reg           irqarray1_soft_re;
wire   [15:0] irqarray1_use_edge;
reg    [15:0] irqarray1_edge_triggered_storage;
reg           irqarray1_edge_triggered_re;
wire   [15:0] irqarray1_rising;
reg    [15:0] irqarray1_polarity_storage;
reg           irqarray1_polarity_re;
wire          irqarray1_eventsourceflex16_status;
reg           irqarray1_eventsourceflex16_pending;
reg           irqarray1_eventsourceflex16_clear;
reg           irqarray1_eventsourceflex16_trigger_d;
reg           irqarray1_eventsourceflex16_trigger_filtered;
wire          irqarray1_eventsourceflex17_status;
reg           irqarray1_eventsourceflex17_pending;
reg           irqarray1_eventsourceflex17_clear;
reg           irqarray1_eventsourceflex17_trigger_d;
reg           irqarray1_eventsourceflex17_trigger_filtered;
wire          irqarray1_eventsourceflex18_status;
reg           irqarray1_eventsourceflex18_pending;
reg           irqarray1_eventsourceflex18_clear;
reg           irqarray1_eventsourceflex18_trigger_d;
reg           irqarray1_eventsourceflex18_trigger_filtered;
wire          irqarray1_eventsourceflex19_status;
reg           irqarray1_eventsourceflex19_pending;
reg           irqarray1_eventsourceflex19_clear;
reg           irqarray1_eventsourceflex19_trigger_d;
reg           irqarray1_eventsourceflex19_trigger_filtered;
wire          irqarray1_eventsourceflex20_status;
reg           irqarray1_eventsourceflex20_pending;
reg           irqarray1_eventsourceflex20_clear;
reg           irqarray1_eventsourceflex20_trigger_d;
reg           irqarray1_eventsourceflex20_trigger_filtered;
wire          irqarray1_eventsourceflex21_status;
reg           irqarray1_eventsourceflex21_pending;
reg           irqarray1_eventsourceflex21_clear;
reg           irqarray1_eventsourceflex21_trigger_d;
reg           irqarray1_eventsourceflex21_trigger_filtered;
wire          irqarray1_eventsourceflex22_status;
reg           irqarray1_eventsourceflex22_pending;
reg           irqarray1_eventsourceflex22_clear;
reg           irqarray1_eventsourceflex22_trigger_d;
reg           irqarray1_eventsourceflex22_trigger_filtered;
wire          irqarray1_eventsourceflex23_status;
reg           irqarray1_eventsourceflex23_pending;
reg           irqarray1_eventsourceflex23_clear;
reg           irqarray1_eventsourceflex23_trigger_d;
reg           irqarray1_eventsourceflex23_trigger_filtered;
wire          irqarray1_eventsourceflex24_status;
reg           irqarray1_eventsourceflex24_pending;
reg           irqarray1_eventsourceflex24_clear;
reg           irqarray1_eventsourceflex24_trigger_d;
reg           irqarray1_eventsourceflex24_trigger_filtered;
wire          irqarray1_eventsourceflex25_status;
reg           irqarray1_eventsourceflex25_pending;
reg           irqarray1_eventsourceflex25_clear;
reg           irqarray1_eventsourceflex25_trigger_d;
reg           irqarray1_eventsourceflex25_trigger_filtered;
wire          irqarray1_eventsourceflex26_status;
reg           irqarray1_eventsourceflex26_pending;
reg           irqarray1_eventsourceflex26_clear;
reg           irqarray1_eventsourceflex26_trigger_d;
reg           irqarray1_eventsourceflex26_trigger_filtered;
wire          irqarray1_eventsourceflex27_status;
reg           irqarray1_eventsourceflex27_pending;
reg           irqarray1_eventsourceflex27_clear;
reg           irqarray1_eventsourceflex27_trigger_d;
reg           irqarray1_eventsourceflex27_trigger_filtered;
wire          irqarray1_eventsourceflex28_status;
reg           irqarray1_eventsourceflex28_pending;
reg           irqarray1_eventsourceflex28_clear;
reg           irqarray1_eventsourceflex28_trigger_d;
reg           irqarray1_eventsourceflex28_trigger_filtered;
wire          irqarray1_eventsourceflex29_status;
reg           irqarray1_eventsourceflex29_pending;
reg           irqarray1_eventsourceflex29_clear;
reg           irqarray1_eventsourceflex29_trigger_d;
reg           irqarray1_eventsourceflex29_trigger_filtered;
wire          irqarray1_eventsourceflex30_status;
reg           irqarray1_eventsourceflex30_pending;
reg           irqarray1_eventsourceflex30_clear;
reg           irqarray1_eventsourceflex30_trigger_d;
reg           irqarray1_eventsourceflex30_trigger_filtered;
wire          irqarray1_eventsourceflex31_status;
reg           irqarray1_eventsourceflex31_pending;
reg           irqarray1_eventsourceflex31_clear;
reg           irqarray1_eventsourceflex31_trigger_d;
reg           irqarray1_eventsourceflex31_trigger_filtered;
wire          irqarray1_usbc_dupe0;
wire          irqarray1_nc_b1s10;
wire          irqarray1_nc_b1s20;
wire          irqarray1_nc_b1s30;
wire          irqarray1_nc_b1s40;
wire          irqarray1_nc_b1s50;
wire          irqarray1_nc_b1s60;
wire          irqarray1_nc_b1s70;
wire          irqarray1_nc_b1s80;
wire          irqarray1_nc_b1s90;
wire          irqarray1_nc_b1s100;
wire          irqarray1_nc_b1s110;
wire          irqarray1_nc_b1s120;
wire          irqarray1_nc_b1s130;
wire          irqarray1_nc_b1s140;
wire          irqarray1_nc_b1s150;
reg    [15:0] irqarray1_status_status;
wire          irqarray1_status_we;
reg           irqarray1_status_re;
wire          irqarray1_usbc_dupe1;
wire          irqarray1_nc_b1s11;
wire          irqarray1_nc_b1s21;
wire          irqarray1_nc_b1s31;
wire          irqarray1_nc_b1s41;
wire          irqarray1_nc_b1s51;
wire          irqarray1_nc_b1s61;
wire          irqarray1_nc_b1s71;
wire          irqarray1_nc_b1s81;
wire          irqarray1_nc_b1s91;
wire          irqarray1_nc_b1s101;
wire          irqarray1_nc_b1s111;
wire          irqarray1_nc_b1s121;
wire          irqarray1_nc_b1s131;
wire          irqarray1_nc_b1s141;
wire          irqarray1_nc_b1s151;
reg    [15:0] irqarray1_pending_status;
wire          irqarray1_pending_we;
reg           irqarray1_pending_re;
reg    [15:0] irqarray1_pending_r;
wire          irqarray1_usbc_dupe2;
wire          irqarray1_nc_b1s12;
wire          irqarray1_nc_b1s22;
wire          irqarray1_nc_b1s32;
wire          irqarray1_nc_b1s42;
wire          irqarray1_nc_b1s52;
wire          irqarray1_nc_b1s62;
wire          irqarray1_nc_b1s72;
wire          irqarray1_nc_b1s82;
wire          irqarray1_nc_b1s92;
wire          irqarray1_nc_b1s102;
wire          irqarray1_nc_b1s112;
wire          irqarray1_nc_b1s122;
wire          irqarray1_nc_b1s132;
wire          irqarray1_nc_b1s142;
wire          irqarray1_nc_b1s152;
reg    [15:0] irqarray1_enable_storage;
reg           irqarray1_enable_re;
wire          irqarray2_irq;
wire   [15:0] irqarray2_interrupts;
reg    [15:0] irqarray2_trigger;
reg    [15:0] irqarray2_soft_storage;
reg           irqarray2_soft_re;
wire   [15:0] irqarray2_use_edge;
reg    [15:0] irqarray2_edge_triggered_storage;
reg           irqarray2_edge_triggered_re;
wire   [15:0] irqarray2_rising;
reg    [15:0] irqarray2_polarity_storage;
reg           irqarray2_polarity_re;
wire          irqarray2_eventsourceflex32_status;
reg           irqarray2_eventsourceflex32_pending;
reg           irqarray2_eventsourceflex32_clear;
reg           irqarray2_eventsourceflex32_trigger_d;
reg           irqarray2_eventsourceflex32_trigger_filtered;
wire          irqarray2_eventsourceflex33_status;
reg           irqarray2_eventsourceflex33_pending;
reg           irqarray2_eventsourceflex33_clear;
reg           irqarray2_eventsourceflex33_trigger_d;
reg           irqarray2_eventsourceflex33_trigger_filtered;
wire          irqarray2_eventsourceflex34_status;
reg           irqarray2_eventsourceflex34_pending;
reg           irqarray2_eventsourceflex34_clear;
reg           irqarray2_eventsourceflex34_trigger_d;
reg           irqarray2_eventsourceflex34_trigger_filtered;
wire          irqarray2_eventsourceflex35_status;
reg           irqarray2_eventsourceflex35_pending;
reg           irqarray2_eventsourceflex35_clear;
reg           irqarray2_eventsourceflex35_trigger_d;
reg           irqarray2_eventsourceflex35_trigger_filtered;
wire          irqarray2_eventsourceflex36_status;
reg           irqarray2_eventsourceflex36_pending;
reg           irqarray2_eventsourceflex36_clear;
reg           irqarray2_eventsourceflex36_trigger_d;
reg           irqarray2_eventsourceflex36_trigger_filtered;
wire          irqarray2_eventsourceflex37_status;
reg           irqarray2_eventsourceflex37_pending;
reg           irqarray2_eventsourceflex37_clear;
reg           irqarray2_eventsourceflex37_trigger_d;
reg           irqarray2_eventsourceflex37_trigger_filtered;
wire          irqarray2_eventsourceflex38_status;
reg           irqarray2_eventsourceflex38_pending;
reg           irqarray2_eventsourceflex38_clear;
reg           irqarray2_eventsourceflex38_trigger_d;
reg           irqarray2_eventsourceflex38_trigger_filtered;
wire          irqarray2_eventsourceflex39_status;
reg           irqarray2_eventsourceflex39_pending;
reg           irqarray2_eventsourceflex39_clear;
reg           irqarray2_eventsourceflex39_trigger_d;
reg           irqarray2_eventsourceflex39_trigger_filtered;
wire          irqarray2_eventsourceflex40_status;
reg           irqarray2_eventsourceflex40_pending;
reg           irqarray2_eventsourceflex40_clear;
reg           irqarray2_eventsourceflex40_trigger_d;
reg           irqarray2_eventsourceflex40_trigger_filtered;
wire          irqarray2_eventsourceflex41_status;
reg           irqarray2_eventsourceflex41_pending;
reg           irqarray2_eventsourceflex41_clear;
reg           irqarray2_eventsourceflex41_trigger_d;
reg           irqarray2_eventsourceflex41_trigger_filtered;
wire          irqarray2_eventsourceflex42_status;
reg           irqarray2_eventsourceflex42_pending;
reg           irqarray2_eventsourceflex42_clear;
reg           irqarray2_eventsourceflex42_trigger_d;
reg           irqarray2_eventsourceflex42_trigger_filtered;
wire          irqarray2_eventsourceflex43_status;
reg           irqarray2_eventsourceflex43_pending;
reg           irqarray2_eventsourceflex43_clear;
reg           irqarray2_eventsourceflex43_trigger_d;
reg           irqarray2_eventsourceflex43_trigger_filtered;
wire          irqarray2_eventsourceflex44_status;
reg           irqarray2_eventsourceflex44_pending;
reg           irqarray2_eventsourceflex44_clear;
reg           irqarray2_eventsourceflex44_trigger_d;
reg           irqarray2_eventsourceflex44_trigger_filtered;
wire          irqarray2_eventsourceflex45_status;
reg           irqarray2_eventsourceflex45_pending;
reg           irqarray2_eventsourceflex45_clear;
reg           irqarray2_eventsourceflex45_trigger_d;
reg           irqarray2_eventsourceflex45_trigger_filtered;
wire          irqarray2_eventsourceflex46_status;
reg           irqarray2_eventsourceflex46_pending;
reg           irqarray2_eventsourceflex46_clear;
reg           irqarray2_eventsourceflex46_trigger_d;
reg           irqarray2_eventsourceflex46_trigger_filtered;
wire          irqarray2_eventsourceflex47_status;
reg           irqarray2_eventsourceflex47_pending;
reg           irqarray2_eventsourceflex47_clear;
reg           irqarray2_eventsourceflex47_trigger_d;
reg           irqarray2_eventsourceflex47_trigger_filtered;
wire          irqarray2_qfcirq0;
wire          irqarray2_mdmairq0;
wire          irqarray2_mbox_irq_available0;
wire          irqarray2_mbox_irq_abort_init0;
wire          irqarray2_mbox_irq_done0;
wire          irqarray2_mbox_irq_error0;
wire          irqarray2_nc_b2s60;
wire          irqarray2_nc_b2s70;
wire          irqarray2_nc_b2s80;
wire          irqarray2_nc_b2s90;
wire          irqarray2_nc_b2s100;
wire          irqarray2_nc_b2s110;
wire          irqarray2_nc_b2s120;
wire          irqarray2_nc_b2s130;
wire          irqarray2_nc_b2s140;
wire          irqarray2_aowkupint0;
reg    [15:0] irqarray2_status_status;
wire          irqarray2_status_we;
reg           irqarray2_status_re;
wire          irqarray2_qfcirq1;
wire          irqarray2_mdmairq1;
wire          irqarray2_mbox_irq_available1;
wire          irqarray2_mbox_irq_abort_init1;
wire          irqarray2_mbox_irq_done1;
wire          irqarray2_mbox_irq_error1;
wire          irqarray2_nc_b2s61;
wire          irqarray2_nc_b2s71;
wire          irqarray2_nc_b2s81;
wire          irqarray2_nc_b2s91;
wire          irqarray2_nc_b2s101;
wire          irqarray2_nc_b2s111;
wire          irqarray2_nc_b2s121;
wire          irqarray2_nc_b2s131;
wire          irqarray2_nc_b2s141;
wire          irqarray2_aowkupint1;
reg    [15:0] irqarray2_pending_status;
wire          irqarray2_pending_we;
reg           irqarray2_pending_re;
reg    [15:0] irqarray2_pending_r;
wire          irqarray2_qfcirq2;
wire          irqarray2_mdmairq2;
wire          irqarray2_mbox_irq_available2;
wire          irqarray2_mbox_irq_abort_init2;
wire          irqarray2_mbox_irq_done2;
wire          irqarray2_mbox_irq_error2;
wire          irqarray2_nc_b2s62;
wire          irqarray2_nc_b2s72;
wire          irqarray2_nc_b2s82;
wire          irqarray2_nc_b2s92;
wire          irqarray2_nc_b2s102;
wire          irqarray2_nc_b2s112;
wire          irqarray2_nc_b2s122;
wire          irqarray2_nc_b2s132;
wire          irqarray2_nc_b2s142;
wire          irqarray2_aowkupint2;
reg    [15:0] irqarray2_enable_storage;
reg           irqarray2_enable_re;
wire          irqarray3_irq;
wire   [15:0] irqarray3_interrupts;
reg    [15:0] irqarray3_trigger;
reg    [15:0] irqarray3_soft_storage;
reg           irqarray3_soft_re;
wire   [15:0] irqarray3_use_edge;
reg    [15:0] irqarray3_edge_triggered_storage;
reg           irqarray3_edge_triggered_re;
wire   [15:0] irqarray3_rising;
reg    [15:0] irqarray3_polarity_storage;
reg           irqarray3_polarity_re;
wire          irqarray3_eventsourceflex48_status;
reg           irqarray3_eventsourceflex48_pending;
reg           irqarray3_eventsourceflex48_clear;
reg           irqarray3_eventsourceflex48_trigger_d;
reg           irqarray3_eventsourceflex48_trigger_filtered;
wire          irqarray3_eventsourceflex49_status;
reg           irqarray3_eventsourceflex49_pending;
reg           irqarray3_eventsourceflex49_clear;
reg           irqarray3_eventsourceflex49_trigger_d;
reg           irqarray3_eventsourceflex49_trigger_filtered;
wire          irqarray3_eventsourceflex50_status;
reg           irqarray3_eventsourceflex50_pending;
reg           irqarray3_eventsourceflex50_clear;
reg           irqarray3_eventsourceflex50_trigger_d;
reg           irqarray3_eventsourceflex50_trigger_filtered;
wire          irqarray3_eventsourceflex51_status;
reg           irqarray3_eventsourceflex51_pending;
reg           irqarray3_eventsourceflex51_clear;
reg           irqarray3_eventsourceflex51_trigger_d;
reg           irqarray3_eventsourceflex51_trigger_filtered;
wire          irqarray3_eventsourceflex52_status;
reg           irqarray3_eventsourceflex52_pending;
reg           irqarray3_eventsourceflex52_clear;
reg           irqarray3_eventsourceflex52_trigger_d;
reg           irqarray3_eventsourceflex52_trigger_filtered;
wire          irqarray3_eventsourceflex53_status;
reg           irqarray3_eventsourceflex53_pending;
reg           irqarray3_eventsourceflex53_clear;
reg           irqarray3_eventsourceflex53_trigger_d;
reg           irqarray3_eventsourceflex53_trigger_filtered;
wire          irqarray3_eventsourceflex54_status;
reg           irqarray3_eventsourceflex54_pending;
reg           irqarray3_eventsourceflex54_clear;
reg           irqarray3_eventsourceflex54_trigger_d;
reg           irqarray3_eventsourceflex54_trigger_filtered;
wire          irqarray3_eventsourceflex55_status;
reg           irqarray3_eventsourceflex55_pending;
reg           irqarray3_eventsourceflex55_clear;
reg           irqarray3_eventsourceflex55_trigger_d;
reg           irqarray3_eventsourceflex55_trigger_filtered;
wire          irqarray3_eventsourceflex56_status;
reg           irqarray3_eventsourceflex56_pending;
reg           irqarray3_eventsourceflex56_clear;
reg           irqarray3_eventsourceflex56_trigger_d;
reg           irqarray3_eventsourceflex56_trigger_filtered;
wire          irqarray3_eventsourceflex57_status;
reg           irqarray3_eventsourceflex57_pending;
reg           irqarray3_eventsourceflex57_clear;
reg           irqarray3_eventsourceflex57_trigger_d;
reg           irqarray3_eventsourceflex57_trigger_filtered;
wire          irqarray3_eventsourceflex58_status;
reg           irqarray3_eventsourceflex58_pending;
reg           irqarray3_eventsourceflex58_clear;
reg           irqarray3_eventsourceflex58_trigger_d;
reg           irqarray3_eventsourceflex58_trigger_filtered;
wire          irqarray3_eventsourceflex59_status;
reg           irqarray3_eventsourceflex59_pending;
reg           irqarray3_eventsourceflex59_clear;
reg           irqarray3_eventsourceflex59_trigger_d;
reg           irqarray3_eventsourceflex59_trigger_filtered;
wire          irqarray3_eventsourceflex60_status;
reg           irqarray3_eventsourceflex60_pending;
reg           irqarray3_eventsourceflex60_clear;
reg           irqarray3_eventsourceflex60_trigger_d;
reg           irqarray3_eventsourceflex60_trigger_filtered;
wire          irqarray3_eventsourceflex61_status;
reg           irqarray3_eventsourceflex61_pending;
reg           irqarray3_eventsourceflex61_clear;
reg           irqarray3_eventsourceflex61_trigger_d;
reg           irqarray3_eventsourceflex61_trigger_filtered;
wire          irqarray3_eventsourceflex62_status;
reg           irqarray3_eventsourceflex62_pending;
reg           irqarray3_eventsourceflex62_clear;
reg           irqarray3_eventsourceflex62_trigger_d;
reg           irqarray3_eventsourceflex62_trigger_filtered;
wire          irqarray3_eventsourceflex63_status;
reg           irqarray3_eventsourceflex63_pending;
reg           irqarray3_eventsourceflex63_clear;
reg           irqarray3_eventsourceflex63_trigger_d;
reg           irqarray3_eventsourceflex63_trigger_filtered;
wire          irqarray3_trng_done0;
wire          irqarray3_aes_done0;
wire          irqarray3_pke_done0;
wire          irqarray3_hash_done0;
wire          irqarray3_alu_done0;
wire          irqarray3_sdma_ichdone0;
wire          irqarray3_sdma_schdone0;
wire          irqarray3_sdma_xchdone0;
wire          irqarray3_nc_b3s80;
wire          irqarray3_nc_b3s90;
wire          irqarray3_nc_b3s100;
wire          irqarray3_nc_b3s110;
wire          irqarray3_nc_b3s120;
wire          irqarray3_nc_b3s130;
wire          irqarray3_nc_b3s140;
wire          irqarray3_nc_b3s150;
reg    [15:0] irqarray3_status_status;
wire          irqarray3_status_we;
reg           irqarray3_status_re;
wire          irqarray3_trng_done1;
wire          irqarray3_aes_done1;
wire          irqarray3_pke_done1;
wire          irqarray3_hash_done1;
wire          irqarray3_alu_done1;
wire          irqarray3_sdma_ichdone1;
wire          irqarray3_sdma_schdone1;
wire          irqarray3_sdma_xchdone1;
wire          irqarray3_nc_b3s81;
wire          irqarray3_nc_b3s91;
wire          irqarray3_nc_b3s101;
wire          irqarray3_nc_b3s111;
wire          irqarray3_nc_b3s121;
wire          irqarray3_nc_b3s131;
wire          irqarray3_nc_b3s141;
wire          irqarray3_nc_b3s151;
reg    [15:0] irqarray3_pending_status;
wire          irqarray3_pending_we;
reg           irqarray3_pending_re;
reg    [15:0] irqarray3_pending_r;
wire          irqarray3_trng_done2;
wire          irqarray3_aes_done2;
wire          irqarray3_pke_done2;
wire          irqarray3_hash_done2;
wire          irqarray3_alu_done2;
wire          irqarray3_sdma_ichdone2;
wire          irqarray3_sdma_schdone2;
wire          irqarray3_sdma_xchdone2;
wire          irqarray3_nc_b3s82;
wire          irqarray3_nc_b3s92;
wire          irqarray3_nc_b3s102;
wire          irqarray3_nc_b3s112;
wire          irqarray3_nc_b3s122;
wire          irqarray3_nc_b3s132;
wire          irqarray3_nc_b3s142;
wire          irqarray3_nc_b3s152;
reg    [15:0] irqarray3_enable_storage;
reg           irqarray3_enable_re;
wire          irqarray4_irq;
wire   [15:0] irqarray4_interrupts;
reg    [15:0] irqarray4_trigger;
reg    [15:0] irqarray4_soft_storage;
reg           irqarray4_soft_re;
wire   [15:0] irqarray4_use_edge;
reg    [15:0] irqarray4_edge_triggered_storage;
reg           irqarray4_edge_triggered_re;
wire   [15:0] irqarray4_rising;
reg    [15:0] irqarray4_polarity_storage;
reg           irqarray4_polarity_re;
wire          irqarray4_eventsourceflex64_status;
reg           irqarray4_eventsourceflex64_pending;
reg           irqarray4_eventsourceflex64_clear;
reg           irqarray4_eventsourceflex64_trigger_d;
reg           irqarray4_eventsourceflex64_trigger_filtered;
wire          irqarray4_eventsourceflex65_status;
reg           irqarray4_eventsourceflex65_pending;
reg           irqarray4_eventsourceflex65_clear;
reg           irqarray4_eventsourceflex65_trigger_d;
reg           irqarray4_eventsourceflex65_trigger_filtered;
wire          irqarray4_eventsourceflex66_status;
reg           irqarray4_eventsourceflex66_pending;
reg           irqarray4_eventsourceflex66_clear;
reg           irqarray4_eventsourceflex66_trigger_d;
reg           irqarray4_eventsourceflex66_trigger_filtered;
wire          irqarray4_eventsourceflex67_status;
reg           irqarray4_eventsourceflex67_pending;
reg           irqarray4_eventsourceflex67_clear;
reg           irqarray4_eventsourceflex67_trigger_d;
reg           irqarray4_eventsourceflex67_trigger_filtered;
wire          irqarray4_eventsourceflex68_status;
reg           irqarray4_eventsourceflex68_pending;
reg           irqarray4_eventsourceflex68_clear;
reg           irqarray4_eventsourceflex68_trigger_d;
reg           irqarray4_eventsourceflex68_trigger_filtered;
wire          irqarray4_eventsourceflex69_status;
reg           irqarray4_eventsourceflex69_pending;
reg           irqarray4_eventsourceflex69_clear;
reg           irqarray4_eventsourceflex69_trigger_d;
reg           irqarray4_eventsourceflex69_trigger_filtered;
wire          irqarray4_eventsourceflex70_status;
reg           irqarray4_eventsourceflex70_pending;
reg           irqarray4_eventsourceflex70_clear;
reg           irqarray4_eventsourceflex70_trigger_d;
reg           irqarray4_eventsourceflex70_trigger_filtered;
wire          irqarray4_eventsourceflex71_status;
reg           irqarray4_eventsourceflex71_pending;
reg           irqarray4_eventsourceflex71_clear;
reg           irqarray4_eventsourceflex71_trigger_d;
reg           irqarray4_eventsourceflex71_trigger_filtered;
wire          irqarray4_eventsourceflex72_status;
reg           irqarray4_eventsourceflex72_pending;
reg           irqarray4_eventsourceflex72_clear;
reg           irqarray4_eventsourceflex72_trigger_d;
reg           irqarray4_eventsourceflex72_trigger_filtered;
wire          irqarray4_eventsourceflex73_status;
reg           irqarray4_eventsourceflex73_pending;
reg           irqarray4_eventsourceflex73_clear;
reg           irqarray4_eventsourceflex73_trigger_d;
reg           irqarray4_eventsourceflex73_trigger_filtered;
wire          irqarray4_eventsourceflex74_status;
reg           irqarray4_eventsourceflex74_pending;
reg           irqarray4_eventsourceflex74_clear;
reg           irqarray4_eventsourceflex74_trigger_d;
reg           irqarray4_eventsourceflex74_trigger_filtered;
wire          irqarray4_eventsourceflex75_status;
reg           irqarray4_eventsourceflex75_pending;
reg           irqarray4_eventsourceflex75_clear;
reg           irqarray4_eventsourceflex75_trigger_d;
reg           irqarray4_eventsourceflex75_trigger_filtered;
wire          irqarray4_eventsourceflex76_status;
reg           irqarray4_eventsourceflex76_pending;
reg           irqarray4_eventsourceflex76_clear;
reg           irqarray4_eventsourceflex76_trigger_d;
reg           irqarray4_eventsourceflex76_trigger_filtered;
wire          irqarray4_eventsourceflex77_status;
reg           irqarray4_eventsourceflex77_pending;
reg           irqarray4_eventsourceflex77_clear;
reg           irqarray4_eventsourceflex77_trigger_d;
reg           irqarray4_eventsourceflex77_trigger_filtered;
wire          irqarray4_eventsourceflex78_status;
reg           irqarray4_eventsourceflex78_pending;
reg           irqarray4_eventsourceflex78_clear;
reg           irqarray4_eventsourceflex78_trigger_d;
reg           irqarray4_eventsourceflex78_trigger_filtered;
wire          irqarray4_eventsourceflex79_status;
reg           irqarray4_eventsourceflex79_pending;
reg           irqarray4_eventsourceflex79_clear;
reg           irqarray4_eventsourceflex79_trigger_d;
reg           irqarray4_eventsourceflex79_trigger_filtered;
wire          irqarray4_trng_done_dupe0;
wire          irqarray4_aes_done_dupe0;
wire          irqarray4_pke_done_dupe0;
wire          irqarray4_hash_done_dupe0;
wire          irqarray4_alu_done_dupe0;
wire          irqarray4_sdma_ichdone_dupe0;
wire          irqarray4_sdma_schdone_dupe0;
wire          irqarray4_sdma_xchdone_dupe0;
wire          irqarray4_nc_b4s80;
wire          irqarray4_nc_b4s90;
wire          irqarray4_nc_b4s100;
wire          irqarray4_nc_b4s110;
wire          irqarray4_nc_b4s120;
wire          irqarray4_nc_b4s130;
wire          irqarray4_nc_b4s140;
wire          irqarray4_nc_b4s150;
reg    [15:0] irqarray4_status_status;
wire          irqarray4_status_we;
reg           irqarray4_status_re;
wire          irqarray4_trng_done_dupe1;
wire          irqarray4_aes_done_dupe1;
wire          irqarray4_pke_done_dupe1;
wire          irqarray4_hash_done_dupe1;
wire          irqarray4_alu_done_dupe1;
wire          irqarray4_sdma_ichdone_dupe1;
wire          irqarray4_sdma_schdone_dupe1;
wire          irqarray4_sdma_xchdone_dupe1;
wire          irqarray4_nc_b4s81;
wire          irqarray4_nc_b4s91;
wire          irqarray4_nc_b4s101;
wire          irqarray4_nc_b4s111;
wire          irqarray4_nc_b4s121;
wire          irqarray4_nc_b4s131;
wire          irqarray4_nc_b4s141;
wire          irqarray4_nc_b4s151;
reg    [15:0] irqarray4_pending_status;
wire          irqarray4_pending_we;
reg           irqarray4_pending_re;
reg    [15:0] irqarray4_pending_r;
wire          irqarray4_trng_done_dupe2;
wire          irqarray4_aes_done_dupe2;
wire          irqarray4_pke_done_dupe2;
wire          irqarray4_hash_done_dupe2;
wire          irqarray4_alu_done_dupe2;
wire          irqarray4_sdma_ichdone_dupe2;
wire          irqarray4_sdma_schdone_dupe2;
wire          irqarray4_sdma_xchdone_dupe2;
wire          irqarray4_nc_b4s82;
wire          irqarray4_nc_b4s92;
wire          irqarray4_nc_b4s102;
wire          irqarray4_nc_b4s112;
wire          irqarray4_nc_b4s122;
wire          irqarray4_nc_b4s132;
wire          irqarray4_nc_b4s142;
wire          irqarray4_nc_b4s152;
reg    [15:0] irqarray4_enable_storage;
reg           irqarray4_enable_re;
wire          irqarray5_irq;
wire   [15:0] irqarray5_interrupts;
reg    [15:0] irqarray5_trigger;
reg    [15:0] irqarray5_soft_storage;
reg           irqarray5_soft_re;
wire   [15:0] irqarray5_use_edge;
reg    [15:0] irqarray5_edge_triggered_storage;
reg           irqarray5_edge_triggered_re;
wire   [15:0] irqarray5_rising;
reg    [15:0] irqarray5_polarity_storage;
reg           irqarray5_polarity_re;
wire          irqarray5_eventsourceflex80_status;
reg           irqarray5_eventsourceflex80_pending;
reg           irqarray5_eventsourceflex80_clear;
reg           irqarray5_eventsourceflex80_trigger_d;
reg           irqarray5_eventsourceflex80_trigger_filtered;
wire          irqarray5_eventsourceflex81_status;
reg           irqarray5_eventsourceflex81_pending;
reg           irqarray5_eventsourceflex81_clear;
reg           irqarray5_eventsourceflex81_trigger_d;
reg           irqarray5_eventsourceflex81_trigger_filtered;
wire          irqarray5_eventsourceflex82_status;
reg           irqarray5_eventsourceflex82_pending;
reg           irqarray5_eventsourceflex82_clear;
reg           irqarray5_eventsourceflex82_trigger_d;
reg           irqarray5_eventsourceflex82_trigger_filtered;
wire          irqarray5_eventsourceflex83_status;
reg           irqarray5_eventsourceflex83_pending;
reg           irqarray5_eventsourceflex83_clear;
reg           irqarray5_eventsourceflex83_trigger_d;
reg           irqarray5_eventsourceflex83_trigger_filtered;
wire          irqarray5_eventsourceflex84_status;
reg           irqarray5_eventsourceflex84_pending;
reg           irqarray5_eventsourceflex84_clear;
reg           irqarray5_eventsourceflex84_trigger_d;
reg           irqarray5_eventsourceflex84_trigger_filtered;
wire          irqarray5_eventsourceflex85_status;
reg           irqarray5_eventsourceflex85_pending;
reg           irqarray5_eventsourceflex85_clear;
reg           irqarray5_eventsourceflex85_trigger_d;
reg           irqarray5_eventsourceflex85_trigger_filtered;
wire          irqarray5_eventsourceflex86_status;
reg           irqarray5_eventsourceflex86_pending;
reg           irqarray5_eventsourceflex86_clear;
reg           irqarray5_eventsourceflex86_trigger_d;
reg           irqarray5_eventsourceflex86_trigger_filtered;
wire          irqarray5_eventsourceflex87_status;
reg           irqarray5_eventsourceflex87_pending;
reg           irqarray5_eventsourceflex87_clear;
reg           irqarray5_eventsourceflex87_trigger_d;
reg           irqarray5_eventsourceflex87_trigger_filtered;
wire          irqarray5_eventsourceflex88_status;
reg           irqarray5_eventsourceflex88_pending;
reg           irqarray5_eventsourceflex88_clear;
reg           irqarray5_eventsourceflex88_trigger_d;
reg           irqarray5_eventsourceflex88_trigger_filtered;
wire          irqarray5_eventsourceflex89_status;
reg           irqarray5_eventsourceflex89_pending;
reg           irqarray5_eventsourceflex89_clear;
reg           irqarray5_eventsourceflex89_trigger_d;
reg           irqarray5_eventsourceflex89_trigger_filtered;
wire          irqarray5_eventsourceflex90_status;
reg           irqarray5_eventsourceflex90_pending;
reg           irqarray5_eventsourceflex90_clear;
reg           irqarray5_eventsourceflex90_trigger_d;
reg           irqarray5_eventsourceflex90_trigger_filtered;
wire          irqarray5_eventsourceflex91_status;
reg           irqarray5_eventsourceflex91_pending;
reg           irqarray5_eventsourceflex91_clear;
reg           irqarray5_eventsourceflex91_trigger_d;
reg           irqarray5_eventsourceflex91_trigger_filtered;
wire          irqarray5_eventsourceflex92_status;
reg           irqarray5_eventsourceflex92_pending;
reg           irqarray5_eventsourceflex92_clear;
reg           irqarray5_eventsourceflex92_trigger_d;
reg           irqarray5_eventsourceflex92_trigger_filtered;
wire          irqarray5_eventsourceflex93_status;
reg           irqarray5_eventsourceflex93_pending;
reg           irqarray5_eventsourceflex93_clear;
reg           irqarray5_eventsourceflex93_trigger_d;
reg           irqarray5_eventsourceflex93_trigger_filtered;
wire          irqarray5_eventsourceflex94_status;
reg           irqarray5_eventsourceflex94_pending;
reg           irqarray5_eventsourceflex94_clear;
reg           irqarray5_eventsourceflex94_trigger_d;
reg           irqarray5_eventsourceflex94_trigger_filtered;
wire          irqarray5_eventsourceflex95_status;
reg           irqarray5_eventsourceflex95_pending;
reg           irqarray5_eventsourceflex95_clear;
reg           irqarray5_eventsourceflex95_trigger_d;
reg           irqarray5_eventsourceflex95_trigger_filtered;
wire          irqarray5_uart0_rx0;
wire          irqarray5_uart0_tx0;
wire          irqarray5_uart0_rx_char0;
wire          irqarray5_uart0_err0;
wire          irqarray5_uart1_rx0;
wire          irqarray5_uart1_tx0;
wire          irqarray5_uart1_rx_char0;
wire          irqarray5_uart1_err0;
wire          irqarray5_uart2_rx0;
wire          irqarray5_uart2_tx0;
wire          irqarray5_uart2_rx_char0;
wire          irqarray5_uart2_err0;
wire          irqarray5_uart3_rx0;
wire          irqarray5_uart3_tx0;
wire          irqarray5_uart3_rx_char0;
wire          irqarray5_uart3_err0;
reg    [15:0] irqarray5_status_status;
wire          irqarray5_status_we;
reg           irqarray5_status_re;
wire          irqarray5_uart0_rx1;
wire          irqarray5_uart0_tx1;
wire          irqarray5_uart0_rx_char1;
wire          irqarray5_uart0_err1;
wire          irqarray5_uart1_rx1;
wire          irqarray5_uart1_tx1;
wire          irqarray5_uart1_rx_char1;
wire          irqarray5_uart1_err1;
wire          irqarray5_uart2_rx1;
wire          irqarray5_uart2_tx1;
wire          irqarray5_uart2_rx_char1;
wire          irqarray5_uart2_err1;
wire          irqarray5_uart3_rx1;
wire          irqarray5_uart3_tx1;
wire          irqarray5_uart3_rx_char1;
wire          irqarray5_uart3_err1;
reg    [15:0] irqarray5_pending_status;
wire          irqarray5_pending_we;
reg           irqarray5_pending_re;
reg    [15:0] irqarray5_pending_r;
wire          irqarray5_uart0_rx2;
wire          irqarray5_uart0_tx2;
wire          irqarray5_uart0_rx_char2;
wire          irqarray5_uart0_err2;
wire          irqarray5_uart1_rx2;
wire          irqarray5_uart1_tx2;
wire          irqarray5_uart1_rx_char2;
wire          irqarray5_uart1_err2;
wire          irqarray5_uart2_rx2;
wire          irqarray5_uart2_tx2;
wire          irqarray5_uart2_rx_char2;
wire          irqarray5_uart2_err2;
wire          irqarray5_uart3_rx2;
wire          irqarray5_uart3_tx2;
wire          irqarray5_uart3_rx_char2;
wire          irqarray5_uart3_err2;
reg    [15:0] irqarray5_enable_storage;
reg           irqarray5_enable_re;
wire          irqarray6_irq;
wire   [15:0] irqarray6_interrupts;
reg    [15:0] irqarray6_trigger;
reg    [15:0] irqarray6_soft_storage;
reg           irqarray6_soft_re;
wire   [15:0] irqarray6_use_edge;
reg    [15:0] irqarray6_edge_triggered_storage;
reg           irqarray6_edge_triggered_re;
wire   [15:0] irqarray6_rising;
reg    [15:0] irqarray6_polarity_storage;
reg           irqarray6_polarity_re;
wire          irqarray6_eventsourceflex96_status;
reg           irqarray6_eventsourceflex96_pending;
reg           irqarray6_eventsourceflex96_clear;
reg           irqarray6_eventsourceflex96_trigger_d;
reg           irqarray6_eventsourceflex96_trigger_filtered;
wire          irqarray6_eventsourceflex97_status;
reg           irqarray6_eventsourceflex97_pending;
reg           irqarray6_eventsourceflex97_clear;
reg           irqarray6_eventsourceflex97_trigger_d;
reg           irqarray6_eventsourceflex97_trigger_filtered;
wire          irqarray6_eventsourceflex98_status;
reg           irqarray6_eventsourceflex98_pending;
reg           irqarray6_eventsourceflex98_clear;
reg           irqarray6_eventsourceflex98_trigger_d;
reg           irqarray6_eventsourceflex98_trigger_filtered;
wire          irqarray6_eventsourceflex99_status;
reg           irqarray6_eventsourceflex99_pending;
reg           irqarray6_eventsourceflex99_clear;
reg           irqarray6_eventsourceflex99_trigger_d;
reg           irqarray6_eventsourceflex99_trigger_filtered;
wire          irqarray6_eventsourceflex100_status;
reg           irqarray6_eventsourceflex100_pending;
reg           irqarray6_eventsourceflex100_clear;
reg           irqarray6_eventsourceflex100_trigger_d;
reg           irqarray6_eventsourceflex100_trigger_filtered;
wire          irqarray6_eventsourceflex101_status;
reg           irqarray6_eventsourceflex101_pending;
reg           irqarray6_eventsourceflex101_clear;
reg           irqarray6_eventsourceflex101_trigger_d;
reg           irqarray6_eventsourceflex101_trigger_filtered;
wire          irqarray6_eventsourceflex102_status;
reg           irqarray6_eventsourceflex102_pending;
reg           irqarray6_eventsourceflex102_clear;
reg           irqarray6_eventsourceflex102_trigger_d;
reg           irqarray6_eventsourceflex102_trigger_filtered;
wire          irqarray6_eventsourceflex103_status;
reg           irqarray6_eventsourceflex103_pending;
reg           irqarray6_eventsourceflex103_clear;
reg           irqarray6_eventsourceflex103_trigger_d;
reg           irqarray6_eventsourceflex103_trigger_filtered;
wire          irqarray6_eventsourceflex104_status;
reg           irqarray6_eventsourceflex104_pending;
reg           irqarray6_eventsourceflex104_clear;
reg           irqarray6_eventsourceflex104_trigger_d;
reg           irqarray6_eventsourceflex104_trigger_filtered;
wire          irqarray6_eventsourceflex105_status;
reg           irqarray6_eventsourceflex105_pending;
reg           irqarray6_eventsourceflex105_clear;
reg           irqarray6_eventsourceflex105_trigger_d;
reg           irqarray6_eventsourceflex105_trigger_filtered;
wire          irqarray6_eventsourceflex106_status;
reg           irqarray6_eventsourceflex106_pending;
reg           irqarray6_eventsourceflex106_clear;
reg           irqarray6_eventsourceflex106_trigger_d;
reg           irqarray6_eventsourceflex106_trigger_filtered;
wire          irqarray6_eventsourceflex107_status;
reg           irqarray6_eventsourceflex107_pending;
reg           irqarray6_eventsourceflex107_clear;
reg           irqarray6_eventsourceflex107_trigger_d;
reg           irqarray6_eventsourceflex107_trigger_filtered;
wire          irqarray6_eventsourceflex108_status;
reg           irqarray6_eventsourceflex108_pending;
reg           irqarray6_eventsourceflex108_clear;
reg           irqarray6_eventsourceflex108_trigger_d;
reg           irqarray6_eventsourceflex108_trigger_filtered;
wire          irqarray6_eventsourceflex109_status;
reg           irqarray6_eventsourceflex109_pending;
reg           irqarray6_eventsourceflex109_clear;
reg           irqarray6_eventsourceflex109_trigger_d;
reg           irqarray6_eventsourceflex109_trigger_filtered;
wire          irqarray6_eventsourceflex110_status;
reg           irqarray6_eventsourceflex110_pending;
reg           irqarray6_eventsourceflex110_clear;
reg           irqarray6_eventsourceflex110_trigger_d;
reg           irqarray6_eventsourceflex110_trigger_filtered;
wire          irqarray6_eventsourceflex111_status;
reg           irqarray6_eventsourceflex111_pending;
reg           irqarray6_eventsourceflex111_clear;
reg           irqarray6_eventsourceflex111_trigger_d;
reg           irqarray6_eventsourceflex111_trigger_filtered;
wire          irqarray6_spim0_rx0;
wire          irqarray6_spim0_tx0;
wire          irqarray6_spim0_cmd0;
wire          irqarray6_spim0_eot0;
wire          irqarray6_spim1_rx0;
wire          irqarray6_spim1_tx0;
wire          irqarray6_spim1_cmd0;
wire          irqarray6_spim1_eot0;
wire          irqarray6_spim2_rx0;
wire          irqarray6_spim2_tx0;
wire          irqarray6_spim2_cmd0;
wire          irqarray6_spim2_eot0;
wire          irqarray6_spim3_rx0;
wire          irqarray6_spim3_tx0;
wire          irqarray6_spim3_cmd0;
wire          irqarray6_spim3_eot0;
reg    [15:0] irqarray6_status_status;
wire          irqarray6_status_we;
reg           irqarray6_status_re;
wire          irqarray6_spim0_rx1;
wire          irqarray6_spim0_tx1;
wire          irqarray6_spim0_cmd1;
wire          irqarray6_spim0_eot1;
wire          irqarray6_spim1_rx1;
wire          irqarray6_spim1_tx1;
wire          irqarray6_spim1_cmd1;
wire          irqarray6_spim1_eot1;
wire          irqarray6_spim2_rx1;
wire          irqarray6_spim2_tx1;
wire          irqarray6_spim2_cmd1;
wire          irqarray6_spim2_eot1;
wire          irqarray6_spim3_rx1;
wire          irqarray6_spim3_tx1;
wire          irqarray6_spim3_cmd1;
wire          irqarray6_spim3_eot1;
reg    [15:0] irqarray6_pending_status;
wire          irqarray6_pending_we;
reg           irqarray6_pending_re;
reg    [15:0] irqarray6_pending_r;
wire          irqarray6_spim0_rx2;
wire          irqarray6_spim0_tx2;
wire          irqarray6_spim0_cmd2;
wire          irqarray6_spim0_eot2;
wire          irqarray6_spim1_rx2;
wire          irqarray6_spim1_tx2;
wire          irqarray6_spim1_cmd2;
wire          irqarray6_spim1_eot2;
wire          irqarray6_spim2_rx2;
wire          irqarray6_spim2_tx2;
wire          irqarray6_spim2_cmd2;
wire          irqarray6_spim2_eot2;
wire          irqarray6_spim3_rx2;
wire          irqarray6_spim3_tx2;
wire          irqarray6_spim3_cmd2;
wire          irqarray6_spim3_eot2;
reg    [15:0] irqarray6_enable_storage;
reg           irqarray6_enable_re;
wire          irqarray7_irq;
wire   [15:0] irqarray7_interrupts;
reg    [15:0] irqarray7_trigger;
reg    [15:0] irqarray7_soft_storage;
reg           irqarray7_soft_re;
wire   [15:0] irqarray7_use_edge;
reg    [15:0] irqarray7_edge_triggered_storage;
reg           irqarray7_edge_triggered_re;
wire   [15:0] irqarray7_rising;
reg    [15:0] irqarray7_polarity_storage;
reg           irqarray7_polarity_re;
wire          irqarray7_eventsourceflex112_status;
reg           irqarray7_eventsourceflex112_pending;
reg           irqarray7_eventsourceflex112_clear;
reg           irqarray7_eventsourceflex112_trigger_d;
reg           irqarray7_eventsourceflex112_trigger_filtered;
wire          irqarray7_eventsourceflex113_status;
reg           irqarray7_eventsourceflex113_pending;
reg           irqarray7_eventsourceflex113_clear;
reg           irqarray7_eventsourceflex113_trigger_d;
reg           irqarray7_eventsourceflex113_trigger_filtered;
wire          irqarray7_eventsourceflex114_status;
reg           irqarray7_eventsourceflex114_pending;
reg           irqarray7_eventsourceflex114_clear;
reg           irqarray7_eventsourceflex114_trigger_d;
reg           irqarray7_eventsourceflex114_trigger_filtered;
wire          irqarray7_eventsourceflex115_status;
reg           irqarray7_eventsourceflex115_pending;
reg           irqarray7_eventsourceflex115_clear;
reg           irqarray7_eventsourceflex115_trigger_d;
reg           irqarray7_eventsourceflex115_trigger_filtered;
wire          irqarray7_eventsourceflex116_status;
reg           irqarray7_eventsourceflex116_pending;
reg           irqarray7_eventsourceflex116_clear;
reg           irqarray7_eventsourceflex116_trigger_d;
reg           irqarray7_eventsourceflex116_trigger_filtered;
wire          irqarray7_eventsourceflex117_status;
reg           irqarray7_eventsourceflex117_pending;
reg           irqarray7_eventsourceflex117_clear;
reg           irqarray7_eventsourceflex117_trigger_d;
reg           irqarray7_eventsourceflex117_trigger_filtered;
wire          irqarray7_eventsourceflex118_status;
reg           irqarray7_eventsourceflex118_pending;
reg           irqarray7_eventsourceflex118_clear;
reg           irqarray7_eventsourceflex118_trigger_d;
reg           irqarray7_eventsourceflex118_trigger_filtered;
wire          irqarray7_eventsourceflex119_status;
reg           irqarray7_eventsourceflex119_pending;
reg           irqarray7_eventsourceflex119_clear;
reg           irqarray7_eventsourceflex119_trigger_d;
reg           irqarray7_eventsourceflex119_trigger_filtered;
wire          irqarray7_eventsourceflex120_status;
reg           irqarray7_eventsourceflex120_pending;
reg           irqarray7_eventsourceflex120_clear;
reg           irqarray7_eventsourceflex120_trigger_d;
reg           irqarray7_eventsourceflex120_trigger_filtered;
wire          irqarray7_eventsourceflex121_status;
reg           irqarray7_eventsourceflex121_pending;
reg           irqarray7_eventsourceflex121_clear;
reg           irqarray7_eventsourceflex121_trigger_d;
reg           irqarray7_eventsourceflex121_trigger_filtered;
wire          irqarray7_eventsourceflex122_status;
reg           irqarray7_eventsourceflex122_pending;
reg           irqarray7_eventsourceflex122_clear;
reg           irqarray7_eventsourceflex122_trigger_d;
reg           irqarray7_eventsourceflex122_trigger_filtered;
wire          irqarray7_eventsourceflex123_status;
reg           irqarray7_eventsourceflex123_pending;
reg           irqarray7_eventsourceflex123_clear;
reg           irqarray7_eventsourceflex123_trigger_d;
reg           irqarray7_eventsourceflex123_trigger_filtered;
wire          irqarray7_eventsourceflex124_status;
reg           irqarray7_eventsourceflex124_pending;
reg           irqarray7_eventsourceflex124_clear;
reg           irqarray7_eventsourceflex124_trigger_d;
reg           irqarray7_eventsourceflex124_trigger_filtered;
wire          irqarray7_eventsourceflex125_status;
reg           irqarray7_eventsourceflex125_pending;
reg           irqarray7_eventsourceflex125_clear;
reg           irqarray7_eventsourceflex125_trigger_d;
reg           irqarray7_eventsourceflex125_trigger_filtered;
wire          irqarray7_eventsourceflex126_status;
reg           irqarray7_eventsourceflex126_pending;
reg           irqarray7_eventsourceflex126_clear;
reg           irqarray7_eventsourceflex126_trigger_d;
reg           irqarray7_eventsourceflex126_trigger_filtered;
wire          irqarray7_eventsourceflex127_status;
reg           irqarray7_eventsourceflex127_pending;
reg           irqarray7_eventsourceflex127_clear;
reg           irqarray7_eventsourceflex127_trigger_d;
reg           irqarray7_eventsourceflex127_trigger_filtered;
wire          irqarray7_i2c0_rx0;
wire          irqarray7_i2c0_tx0;
wire          irqarray7_i2c0_cmd0;
wire          irqarray7_i2c0_eot0;
wire          irqarray7_i2c1_rx0;
wire          irqarray7_i2c1_tx0;
wire          irqarray7_i2c1_cmd0;
wire          irqarray7_i2c1_eot0;
wire          irqarray7_i2c2_rx0;
wire          irqarray7_i2c2_tx0;
wire          irqarray7_i2c2_cmd0;
wire          irqarray7_i2c2_eot0;
wire          irqarray7_i2c3_rx0;
wire          irqarray7_i2c3_tx0;
wire          irqarray7_i2c3_cmd0;
wire          irqarray7_i2c3_eot0;
reg    [15:0] irqarray7_status_status;
wire          irqarray7_status_we;
reg           irqarray7_status_re;
wire          irqarray7_i2c0_rx1;
wire          irqarray7_i2c0_tx1;
wire          irqarray7_i2c0_cmd1;
wire          irqarray7_i2c0_eot1;
wire          irqarray7_i2c1_rx1;
wire          irqarray7_i2c1_tx1;
wire          irqarray7_i2c1_cmd1;
wire          irqarray7_i2c1_eot1;
wire          irqarray7_i2c2_rx1;
wire          irqarray7_i2c2_tx1;
wire          irqarray7_i2c2_cmd1;
wire          irqarray7_i2c2_eot1;
wire          irqarray7_i2c3_rx1;
wire          irqarray7_i2c3_tx1;
wire          irqarray7_i2c3_cmd1;
wire          irqarray7_i2c3_eot1;
reg    [15:0] irqarray7_pending_status;
wire          irqarray7_pending_we;
reg           irqarray7_pending_re;
reg    [15:0] irqarray7_pending_r;
wire          irqarray7_i2c0_rx2;
wire          irqarray7_i2c0_tx2;
wire          irqarray7_i2c0_cmd2;
wire          irqarray7_i2c0_eot2;
wire          irqarray7_i2c1_rx2;
wire          irqarray7_i2c1_tx2;
wire          irqarray7_i2c1_cmd2;
wire          irqarray7_i2c1_eot2;
wire          irqarray7_i2c2_rx2;
wire          irqarray7_i2c2_tx2;
wire          irqarray7_i2c2_cmd2;
wire          irqarray7_i2c2_eot2;
wire          irqarray7_i2c3_rx2;
wire          irqarray7_i2c3_tx2;
wire          irqarray7_i2c3_cmd2;
wire          irqarray7_i2c3_eot2;
reg    [15:0] irqarray7_enable_storage;
reg           irqarray7_enable_re;
wire          irqarray8_irq;
wire   [15:0] irqarray8_interrupts;
reg    [15:0] irqarray8_trigger;
reg    [15:0] irqarray8_soft_storage;
reg           irqarray8_soft_re;
wire   [15:0] irqarray8_use_edge;
reg    [15:0] irqarray8_edge_triggered_storage;
reg           irqarray8_edge_triggered_re;
wire   [15:0] irqarray8_rising;
reg    [15:0] irqarray8_polarity_storage;
reg           irqarray8_polarity_re;
wire          irqarray8_eventsourceflex128_status;
reg           irqarray8_eventsourceflex128_pending;
reg           irqarray8_eventsourceflex128_clear;
reg           irqarray8_eventsourceflex128_trigger_d;
reg           irqarray8_eventsourceflex128_trigger_filtered;
wire          irqarray8_eventsourceflex129_status;
reg           irqarray8_eventsourceflex129_pending;
reg           irqarray8_eventsourceflex129_clear;
reg           irqarray8_eventsourceflex129_trigger_d;
reg           irqarray8_eventsourceflex129_trigger_filtered;
wire          irqarray8_eventsourceflex130_status;
reg           irqarray8_eventsourceflex130_pending;
reg           irqarray8_eventsourceflex130_clear;
reg           irqarray8_eventsourceflex130_trigger_d;
reg           irqarray8_eventsourceflex130_trigger_filtered;
wire          irqarray8_eventsourceflex131_status;
reg           irqarray8_eventsourceflex131_pending;
reg           irqarray8_eventsourceflex131_clear;
reg           irqarray8_eventsourceflex131_trigger_d;
reg           irqarray8_eventsourceflex131_trigger_filtered;
wire          irqarray8_eventsourceflex132_status;
reg           irqarray8_eventsourceflex132_pending;
reg           irqarray8_eventsourceflex132_clear;
reg           irqarray8_eventsourceflex132_trigger_d;
reg           irqarray8_eventsourceflex132_trigger_filtered;
wire          irqarray8_eventsourceflex133_status;
reg           irqarray8_eventsourceflex133_pending;
reg           irqarray8_eventsourceflex133_clear;
reg           irqarray8_eventsourceflex133_trigger_d;
reg           irqarray8_eventsourceflex133_trigger_filtered;
wire          irqarray8_eventsourceflex134_status;
reg           irqarray8_eventsourceflex134_pending;
reg           irqarray8_eventsourceflex134_clear;
reg           irqarray8_eventsourceflex134_trigger_d;
reg           irqarray8_eventsourceflex134_trigger_filtered;
wire          irqarray8_eventsourceflex135_status;
reg           irqarray8_eventsourceflex135_pending;
reg           irqarray8_eventsourceflex135_clear;
reg           irqarray8_eventsourceflex135_trigger_d;
reg           irqarray8_eventsourceflex135_trigger_filtered;
wire          irqarray8_eventsourceflex136_status;
reg           irqarray8_eventsourceflex136_pending;
reg           irqarray8_eventsourceflex136_clear;
reg           irqarray8_eventsourceflex136_trigger_d;
reg           irqarray8_eventsourceflex136_trigger_filtered;
wire          irqarray8_eventsourceflex137_status;
reg           irqarray8_eventsourceflex137_pending;
reg           irqarray8_eventsourceflex137_clear;
reg           irqarray8_eventsourceflex137_trigger_d;
reg           irqarray8_eventsourceflex137_trigger_filtered;
wire          irqarray8_eventsourceflex138_status;
reg           irqarray8_eventsourceflex138_pending;
reg           irqarray8_eventsourceflex138_clear;
reg           irqarray8_eventsourceflex138_trigger_d;
reg           irqarray8_eventsourceflex138_trigger_filtered;
wire          irqarray8_eventsourceflex139_status;
reg           irqarray8_eventsourceflex139_pending;
reg           irqarray8_eventsourceflex139_clear;
reg           irqarray8_eventsourceflex139_trigger_d;
reg           irqarray8_eventsourceflex139_trigger_filtered;
wire          irqarray8_eventsourceflex140_status;
reg           irqarray8_eventsourceflex140_pending;
reg           irqarray8_eventsourceflex140_clear;
reg           irqarray8_eventsourceflex140_trigger_d;
reg           irqarray8_eventsourceflex140_trigger_filtered;
wire          irqarray8_eventsourceflex141_status;
reg           irqarray8_eventsourceflex141_pending;
reg           irqarray8_eventsourceflex141_clear;
reg           irqarray8_eventsourceflex141_trigger_d;
reg           irqarray8_eventsourceflex141_trigger_filtered;
wire          irqarray8_eventsourceflex142_status;
reg           irqarray8_eventsourceflex142_pending;
reg           irqarray8_eventsourceflex142_clear;
reg           irqarray8_eventsourceflex142_trigger_d;
reg           irqarray8_eventsourceflex142_trigger_filtered;
wire          irqarray8_eventsourceflex143_status;
reg           irqarray8_eventsourceflex143_pending;
reg           irqarray8_eventsourceflex143_clear;
reg           irqarray8_eventsourceflex143_trigger_d;
reg           irqarray8_eventsourceflex143_trigger_filtered;
wire          irqarray8_sdio_rx0;
wire          irqarray8_sdio_tx0;
wire          irqarray8_sdio_eot0;
wire          irqarray8_sdio_err0;
wire          irqarray8_i2s_rx0;
wire          irqarray8_i2s_tx0;
wire          irqarray8_nc_b8s60;
wire          irqarray8_nc_b8s70;
wire          irqarray8_cam_rx0;
wire          irqarray8_adc_rx0;
wire          irqarray8_nc_b8s100;
wire          irqarray8_nc_b8s110;
wire          irqarray8_filter_eot0;
wire          irqarray8_filter_act0;
wire          irqarray8_nc_b8s140;
wire          irqarray8_nc_b8s150;
reg    [15:0] irqarray8_status_status;
wire          irqarray8_status_we;
reg           irqarray8_status_re;
wire          irqarray8_sdio_rx1;
wire          irqarray8_sdio_tx1;
wire          irqarray8_sdio_eot1;
wire          irqarray8_sdio_err1;
wire          irqarray8_i2s_rx1;
wire          irqarray8_i2s_tx1;
wire          irqarray8_nc_b8s61;
wire          irqarray8_nc_b8s71;
wire          irqarray8_cam_rx1;
wire          irqarray8_adc_rx1;
wire          irqarray8_nc_b8s101;
wire          irqarray8_nc_b8s111;
wire          irqarray8_filter_eot1;
wire          irqarray8_filter_act1;
wire          irqarray8_nc_b8s141;
wire          irqarray8_nc_b8s151;
reg    [15:0] irqarray8_pending_status;
wire          irqarray8_pending_we;
reg           irqarray8_pending_re;
reg    [15:0] irqarray8_pending_r;
wire          irqarray8_sdio_rx2;
wire          irqarray8_sdio_tx2;
wire          irqarray8_sdio_eot2;
wire          irqarray8_sdio_err2;
wire          irqarray8_i2s_rx2;
wire          irqarray8_i2s_tx2;
wire          irqarray8_nc_b8s62;
wire          irqarray8_nc_b8s72;
wire          irqarray8_cam_rx2;
wire          irqarray8_adc_rx2;
wire          irqarray8_nc_b8s102;
wire          irqarray8_nc_b8s112;
wire          irqarray8_filter_eot2;
wire          irqarray8_filter_act2;
wire          irqarray8_nc_b8s142;
wire          irqarray8_nc_b8s152;
reg    [15:0] irqarray8_enable_storage;
reg           irqarray8_enable_re;
wire          irqarray9_irq;
wire   [15:0] irqarray9_interrupts;
reg    [15:0] irqarray9_trigger;
reg    [15:0] irqarray9_soft_storage;
reg           irqarray9_soft_re;
wire   [15:0] irqarray9_use_edge;
reg    [15:0] irqarray9_edge_triggered_storage;
reg           irqarray9_edge_triggered_re;
wire   [15:0] irqarray9_rising;
reg    [15:0] irqarray9_polarity_storage;
reg           irqarray9_polarity_re;
wire          irqarray9_eventsourceflex144_status;
reg           irqarray9_eventsourceflex144_pending;
reg           irqarray9_eventsourceflex144_clear;
reg           irqarray9_eventsourceflex144_trigger_d;
reg           irqarray9_eventsourceflex144_trigger_filtered;
wire          irqarray9_eventsourceflex145_status;
reg           irqarray9_eventsourceflex145_pending;
reg           irqarray9_eventsourceflex145_clear;
reg           irqarray9_eventsourceflex145_trigger_d;
reg           irqarray9_eventsourceflex145_trigger_filtered;
wire          irqarray9_eventsourceflex146_status;
reg           irqarray9_eventsourceflex146_pending;
reg           irqarray9_eventsourceflex146_clear;
reg           irqarray9_eventsourceflex146_trigger_d;
reg           irqarray9_eventsourceflex146_trigger_filtered;
wire          irqarray9_eventsourceflex147_status;
reg           irqarray9_eventsourceflex147_pending;
reg           irqarray9_eventsourceflex147_clear;
reg           irqarray9_eventsourceflex147_trigger_d;
reg           irqarray9_eventsourceflex147_trigger_filtered;
wire          irqarray9_eventsourceflex148_status;
reg           irqarray9_eventsourceflex148_pending;
reg           irqarray9_eventsourceflex148_clear;
reg           irqarray9_eventsourceflex148_trigger_d;
reg           irqarray9_eventsourceflex148_trigger_filtered;
wire          irqarray9_eventsourceflex149_status;
reg           irqarray9_eventsourceflex149_pending;
reg           irqarray9_eventsourceflex149_clear;
reg           irqarray9_eventsourceflex149_trigger_d;
reg           irqarray9_eventsourceflex149_trigger_filtered;
wire          irqarray9_eventsourceflex150_status;
reg           irqarray9_eventsourceflex150_pending;
reg           irqarray9_eventsourceflex150_clear;
reg           irqarray9_eventsourceflex150_trigger_d;
reg           irqarray9_eventsourceflex150_trigger_filtered;
wire          irqarray9_eventsourceflex151_status;
reg           irqarray9_eventsourceflex151_pending;
reg           irqarray9_eventsourceflex151_clear;
reg           irqarray9_eventsourceflex151_trigger_d;
reg           irqarray9_eventsourceflex151_trigger_filtered;
wire          irqarray9_eventsourceflex152_status;
reg           irqarray9_eventsourceflex152_pending;
reg           irqarray9_eventsourceflex152_clear;
reg           irqarray9_eventsourceflex152_trigger_d;
reg           irqarray9_eventsourceflex152_trigger_filtered;
wire          irqarray9_eventsourceflex153_status;
reg           irqarray9_eventsourceflex153_pending;
reg           irqarray9_eventsourceflex153_clear;
reg           irqarray9_eventsourceflex153_trigger_d;
reg           irqarray9_eventsourceflex153_trigger_filtered;
wire          irqarray9_eventsourceflex154_status;
reg           irqarray9_eventsourceflex154_pending;
reg           irqarray9_eventsourceflex154_clear;
reg           irqarray9_eventsourceflex154_trigger_d;
reg           irqarray9_eventsourceflex154_trigger_filtered;
wire          irqarray9_eventsourceflex155_status;
reg           irqarray9_eventsourceflex155_pending;
reg           irqarray9_eventsourceflex155_clear;
reg           irqarray9_eventsourceflex155_trigger_d;
reg           irqarray9_eventsourceflex155_trigger_filtered;
wire          irqarray9_eventsourceflex156_status;
reg           irqarray9_eventsourceflex156_pending;
reg           irqarray9_eventsourceflex156_clear;
reg           irqarray9_eventsourceflex156_trigger_d;
reg           irqarray9_eventsourceflex156_trigger_filtered;
wire          irqarray9_eventsourceflex157_status;
reg           irqarray9_eventsourceflex157_pending;
reg           irqarray9_eventsourceflex157_clear;
reg           irqarray9_eventsourceflex157_trigger_d;
reg           irqarray9_eventsourceflex157_trigger_filtered;
wire          irqarray9_eventsourceflex158_status;
reg           irqarray9_eventsourceflex158_pending;
reg           irqarray9_eventsourceflex158_clear;
reg           irqarray9_eventsourceflex158_trigger_d;
reg           irqarray9_eventsourceflex158_trigger_filtered;
wire          irqarray9_eventsourceflex159_status;
reg           irqarray9_eventsourceflex159_pending;
reg           irqarray9_eventsourceflex159_clear;
reg           irqarray9_eventsourceflex159_trigger_d;
reg           irqarray9_eventsourceflex159_trigger_filtered;
wire          irqarray9_scif_rx0;
wire          irqarray9_scif_tx0;
wire          irqarray9_scif_rx_char0;
wire          irqarray9_scif_err0;
wire          irqarray9_spis0_rx0;
wire          irqarray9_spis0_tx0;
wire          irqarray9_spis0_eot0;
wire          irqarray9_nc_b9s70;
wire          irqarray9_spis1_rx0;
wire          irqarray9_spis1_tx0;
wire          irqarray9_spis1_eot0;
wire          irqarray9_nc_b9s110;
wire          irqarray9_pwm0_ev0;
wire          irqarray9_pwm1_ev0;
wire          irqarray9_pwm2_ev0;
wire          irqarray9_pwm3_ev0;
reg    [15:0] irqarray9_status_status;
wire          irqarray9_status_we;
reg           irqarray9_status_re;
wire          irqarray9_scif_rx1;
wire          irqarray9_scif_tx1;
wire          irqarray9_scif_rx_char1;
wire          irqarray9_scif_err1;
wire          irqarray9_spis0_rx1;
wire          irqarray9_spis0_tx1;
wire          irqarray9_spis0_eot1;
wire          irqarray9_nc_b9s71;
wire          irqarray9_spis1_rx1;
wire          irqarray9_spis1_tx1;
wire          irqarray9_spis1_eot1;
wire          irqarray9_nc_b9s111;
wire          irqarray9_pwm0_ev1;
wire          irqarray9_pwm1_ev1;
wire          irqarray9_pwm2_ev1;
wire          irqarray9_pwm3_ev1;
reg    [15:0] irqarray9_pending_status;
wire          irqarray9_pending_we;
reg           irqarray9_pending_re;
reg    [15:0] irqarray9_pending_r;
wire          irqarray9_scif_rx2;
wire          irqarray9_scif_tx2;
wire          irqarray9_scif_rx_char2;
wire          irqarray9_scif_err2;
wire          irqarray9_spis0_rx2;
wire          irqarray9_spis0_tx2;
wire          irqarray9_spis0_eot2;
wire          irqarray9_nc_b9s72;
wire          irqarray9_spis1_rx2;
wire          irqarray9_spis1_tx2;
wire          irqarray9_spis1_eot2;
wire          irqarray9_nc_b9s112;
wire          irqarray9_pwm0_ev2;
wire          irqarray9_pwm1_ev2;
wire          irqarray9_pwm2_ev2;
wire          irqarray9_pwm3_ev2;
reg    [15:0] irqarray9_enable_storage;
reg           irqarray9_enable_re;
wire          irqarray10_irq;
wire   [15:0] irqarray10_interrupts;
reg    [15:0] irqarray10_trigger;
reg    [15:0] irqarray10_soft_storage;
reg           irqarray10_soft_re;
wire   [15:0] irqarray10_use_edge;
reg    [15:0] irqarray10_edge_triggered_storage;
reg           irqarray10_edge_triggered_re;
wire   [15:0] irqarray10_rising;
reg    [15:0] irqarray10_polarity_storage;
reg           irqarray10_polarity_re;
wire          irqarray10_eventsourceflex160_status;
reg           irqarray10_eventsourceflex160_pending;
reg           irqarray10_eventsourceflex160_clear;
reg           irqarray10_eventsourceflex160_trigger_d;
reg           irqarray10_eventsourceflex160_trigger_filtered;
wire          irqarray10_eventsourceflex161_status;
reg           irqarray10_eventsourceflex161_pending;
reg           irqarray10_eventsourceflex161_clear;
reg           irqarray10_eventsourceflex161_trigger_d;
reg           irqarray10_eventsourceflex161_trigger_filtered;
wire          irqarray10_eventsourceflex162_status;
reg           irqarray10_eventsourceflex162_pending;
reg           irqarray10_eventsourceflex162_clear;
reg           irqarray10_eventsourceflex162_trigger_d;
reg           irqarray10_eventsourceflex162_trigger_filtered;
wire          irqarray10_eventsourceflex163_status;
reg           irqarray10_eventsourceflex163_pending;
reg           irqarray10_eventsourceflex163_clear;
reg           irqarray10_eventsourceflex163_trigger_d;
reg           irqarray10_eventsourceflex163_trigger_filtered;
wire          irqarray10_eventsourceflex164_status;
reg           irqarray10_eventsourceflex164_pending;
reg           irqarray10_eventsourceflex164_clear;
reg           irqarray10_eventsourceflex164_trigger_d;
reg           irqarray10_eventsourceflex164_trigger_filtered;
wire          irqarray10_eventsourceflex165_status;
reg           irqarray10_eventsourceflex165_pending;
reg           irqarray10_eventsourceflex165_clear;
reg           irqarray10_eventsourceflex165_trigger_d;
reg           irqarray10_eventsourceflex165_trigger_filtered;
wire          irqarray10_eventsourceflex166_status;
reg           irqarray10_eventsourceflex166_pending;
reg           irqarray10_eventsourceflex166_clear;
reg           irqarray10_eventsourceflex166_trigger_d;
reg           irqarray10_eventsourceflex166_trigger_filtered;
wire          irqarray10_eventsourceflex167_status;
reg           irqarray10_eventsourceflex167_pending;
reg           irqarray10_eventsourceflex167_clear;
reg           irqarray10_eventsourceflex167_trigger_d;
reg           irqarray10_eventsourceflex167_trigger_filtered;
wire          irqarray10_eventsourceflex168_status;
reg           irqarray10_eventsourceflex168_pending;
reg           irqarray10_eventsourceflex168_clear;
reg           irqarray10_eventsourceflex168_trigger_d;
reg           irqarray10_eventsourceflex168_trigger_filtered;
wire          irqarray10_eventsourceflex169_status;
reg           irqarray10_eventsourceflex169_pending;
reg           irqarray10_eventsourceflex169_clear;
reg           irqarray10_eventsourceflex169_trigger_d;
reg           irqarray10_eventsourceflex169_trigger_filtered;
wire          irqarray10_eventsourceflex170_status;
reg           irqarray10_eventsourceflex170_pending;
reg           irqarray10_eventsourceflex170_clear;
reg           irqarray10_eventsourceflex170_trigger_d;
reg           irqarray10_eventsourceflex170_trigger_filtered;
wire          irqarray10_eventsourceflex171_status;
reg           irqarray10_eventsourceflex171_pending;
reg           irqarray10_eventsourceflex171_clear;
reg           irqarray10_eventsourceflex171_trigger_d;
reg           irqarray10_eventsourceflex171_trigger_filtered;
wire          irqarray10_eventsourceflex172_status;
reg           irqarray10_eventsourceflex172_pending;
reg           irqarray10_eventsourceflex172_clear;
reg           irqarray10_eventsourceflex172_trigger_d;
reg           irqarray10_eventsourceflex172_trigger_filtered;
wire          irqarray10_eventsourceflex173_status;
reg           irqarray10_eventsourceflex173_pending;
reg           irqarray10_eventsourceflex173_clear;
reg           irqarray10_eventsourceflex173_trigger_d;
reg           irqarray10_eventsourceflex173_trigger_filtered;
wire          irqarray10_eventsourceflex174_status;
reg           irqarray10_eventsourceflex174_pending;
reg           irqarray10_eventsourceflex174_clear;
reg           irqarray10_eventsourceflex174_trigger_d;
reg           irqarray10_eventsourceflex174_trigger_filtered;
wire          irqarray10_eventsourceflex175_status;
reg           irqarray10_eventsourceflex175_pending;
reg           irqarray10_eventsourceflex175_clear;
reg           irqarray10_eventsourceflex175_trigger_d;
reg           irqarray10_eventsourceflex175_trigger_filtered;
wire          irqarray10_ioxirq0;
wire          irqarray10_usbc0;
wire          irqarray10_sddcirq0;
wire          irqarray10_pioirq00;
wire          irqarray10_pioirq10;
wire          irqarray10_pioirq20;
wire          irqarray10_pioirq30;
wire          irqarray10_nc_b10s70;
wire          irqarray10_nc_b10s80;
wire          irqarray10_nc_b10s90;
wire          irqarray10_nc_b10s100;
wire          irqarray10_nc_b10s110;
wire          irqarray10_nc_b10s120;
wire          irqarray10_nc_b10s130;
wire          irqarray10_nc_b10s140;
wire          irqarray10_nc_b10s150;
reg    [15:0] irqarray10_status_status;
wire          irqarray10_status_we;
reg           irqarray10_status_re;
wire          irqarray10_ioxirq1;
wire          irqarray10_usbc1;
wire          irqarray10_sddcirq1;
wire          irqarray10_pioirq01;
wire          irqarray10_pioirq11;
wire          irqarray10_pioirq21;
wire          irqarray10_pioirq31;
wire          irqarray10_nc_b10s71;
wire          irqarray10_nc_b10s81;
wire          irqarray10_nc_b10s91;
wire          irqarray10_nc_b10s101;
wire          irqarray10_nc_b10s111;
wire          irqarray10_nc_b10s121;
wire          irqarray10_nc_b10s131;
wire          irqarray10_nc_b10s141;
wire          irqarray10_nc_b10s151;
reg    [15:0] irqarray10_pending_status;
wire          irqarray10_pending_we;
reg           irqarray10_pending_re;
reg    [15:0] irqarray10_pending_r;
wire          irqarray10_ioxirq2;
wire          irqarray10_usbc2;
wire          irqarray10_sddcirq2;
wire          irqarray10_pioirq02;
wire          irqarray10_pioirq12;
wire          irqarray10_pioirq22;
wire          irqarray10_pioirq32;
wire          irqarray10_nc_b10s72;
wire          irqarray10_nc_b10s82;
wire          irqarray10_nc_b10s92;
wire          irqarray10_nc_b10s102;
wire          irqarray10_nc_b10s112;
wire          irqarray10_nc_b10s122;
wire          irqarray10_nc_b10s132;
wire          irqarray10_nc_b10s142;
wire          irqarray10_nc_b10s152;
reg    [15:0] irqarray10_enable_storage;
reg           irqarray10_enable_re;
wire          irqarray11_irq;
wire   [15:0] irqarray11_interrupts;
reg    [15:0] irqarray11_trigger;
reg    [15:0] irqarray11_soft_storage;
reg           irqarray11_soft_re;
wire   [15:0] irqarray11_use_edge;
reg    [15:0] irqarray11_edge_triggered_storage;
reg           irqarray11_edge_triggered_re;
wire   [15:0] irqarray11_rising;
reg    [15:0] irqarray11_polarity_storage;
reg           irqarray11_polarity_re;
wire          irqarray11_eventsourceflex176_status;
reg           irqarray11_eventsourceflex176_pending;
reg           irqarray11_eventsourceflex176_clear;
reg           irqarray11_eventsourceflex176_trigger_d;
reg           irqarray11_eventsourceflex176_trigger_filtered;
wire          irqarray11_eventsourceflex177_status;
reg           irqarray11_eventsourceflex177_pending;
reg           irqarray11_eventsourceflex177_clear;
reg           irqarray11_eventsourceflex177_trigger_d;
reg           irqarray11_eventsourceflex177_trigger_filtered;
wire          irqarray11_eventsourceflex178_status;
reg           irqarray11_eventsourceflex178_pending;
reg           irqarray11_eventsourceflex178_clear;
reg           irqarray11_eventsourceflex178_trigger_d;
reg           irqarray11_eventsourceflex178_trigger_filtered;
wire          irqarray11_eventsourceflex179_status;
reg           irqarray11_eventsourceflex179_pending;
reg           irqarray11_eventsourceflex179_clear;
reg           irqarray11_eventsourceflex179_trigger_d;
reg           irqarray11_eventsourceflex179_trigger_filtered;
wire          irqarray11_eventsourceflex180_status;
reg           irqarray11_eventsourceflex180_pending;
reg           irqarray11_eventsourceflex180_clear;
reg           irqarray11_eventsourceflex180_trigger_d;
reg           irqarray11_eventsourceflex180_trigger_filtered;
wire          irqarray11_eventsourceflex181_status;
reg           irqarray11_eventsourceflex181_pending;
reg           irqarray11_eventsourceflex181_clear;
reg           irqarray11_eventsourceflex181_trigger_d;
reg           irqarray11_eventsourceflex181_trigger_filtered;
wire          irqarray11_eventsourceflex182_status;
reg           irqarray11_eventsourceflex182_pending;
reg           irqarray11_eventsourceflex182_clear;
reg           irqarray11_eventsourceflex182_trigger_d;
reg           irqarray11_eventsourceflex182_trigger_filtered;
wire          irqarray11_eventsourceflex183_status;
reg           irqarray11_eventsourceflex183_pending;
reg           irqarray11_eventsourceflex183_clear;
reg           irqarray11_eventsourceflex183_trigger_d;
reg           irqarray11_eventsourceflex183_trigger_filtered;
wire          irqarray11_eventsourceflex184_status;
reg           irqarray11_eventsourceflex184_pending;
reg           irqarray11_eventsourceflex184_clear;
reg           irqarray11_eventsourceflex184_trigger_d;
reg           irqarray11_eventsourceflex184_trigger_filtered;
wire          irqarray11_eventsourceflex185_status;
reg           irqarray11_eventsourceflex185_pending;
reg           irqarray11_eventsourceflex185_clear;
reg           irqarray11_eventsourceflex185_trigger_d;
reg           irqarray11_eventsourceflex185_trigger_filtered;
wire          irqarray11_eventsourceflex186_status;
reg           irqarray11_eventsourceflex186_pending;
reg           irqarray11_eventsourceflex186_clear;
reg           irqarray11_eventsourceflex186_trigger_d;
reg           irqarray11_eventsourceflex186_trigger_filtered;
wire          irqarray11_eventsourceflex187_status;
reg           irqarray11_eventsourceflex187_pending;
reg           irqarray11_eventsourceflex187_clear;
reg           irqarray11_eventsourceflex187_trigger_d;
reg           irqarray11_eventsourceflex187_trigger_filtered;
wire          irqarray11_eventsourceflex188_status;
reg           irqarray11_eventsourceflex188_pending;
reg           irqarray11_eventsourceflex188_clear;
reg           irqarray11_eventsourceflex188_trigger_d;
reg           irqarray11_eventsourceflex188_trigger_filtered;
wire          irqarray11_eventsourceflex189_status;
reg           irqarray11_eventsourceflex189_pending;
reg           irqarray11_eventsourceflex189_clear;
reg           irqarray11_eventsourceflex189_trigger_d;
reg           irqarray11_eventsourceflex189_trigger_filtered;
wire          irqarray11_eventsourceflex190_status;
reg           irqarray11_eventsourceflex190_pending;
reg           irqarray11_eventsourceflex190_clear;
reg           irqarray11_eventsourceflex190_trigger_d;
reg           irqarray11_eventsourceflex190_trigger_filtered;
wire          irqarray11_eventsourceflex191_status;
reg           irqarray11_eventsourceflex191_pending;
reg           irqarray11_eventsourceflex191_clear;
reg           irqarray11_eventsourceflex191_trigger_d;
reg           irqarray11_eventsourceflex191_trigger_filtered;
wire          irqarray11_i2s_rx_dupe0;
wire          irqarray11_i2s_tx_dupe0;
wire          irqarray11_nc_b11s20;
wire          irqarray11_nc_b11s30;
wire          irqarray11_nc_b11s40;
wire          irqarray11_nc_b11s50;
wire          irqarray11_nc_b11s60;
wire          irqarray11_nc_b11s70;
wire          irqarray11_nc_b11s80;
wire          irqarray11_nc_b11s90;
wire          irqarray11_nc_b11s100;
wire          irqarray11_nc_b11s110;
wire          irqarray11_nc_b11s120;
wire          irqarray11_nc_b11s130;
wire          irqarray11_nc_b11s140;
wire          irqarray11_nc_b11s150;
reg    [15:0] irqarray11_status_status;
wire          irqarray11_status_we;
reg           irqarray11_status_re;
wire          irqarray11_i2s_rx_dupe1;
wire          irqarray11_i2s_tx_dupe1;
wire          irqarray11_nc_b11s21;
wire          irqarray11_nc_b11s31;
wire          irqarray11_nc_b11s41;
wire          irqarray11_nc_b11s51;
wire          irqarray11_nc_b11s61;
wire          irqarray11_nc_b11s71;
wire          irqarray11_nc_b11s81;
wire          irqarray11_nc_b11s91;
wire          irqarray11_nc_b11s101;
wire          irqarray11_nc_b11s111;
wire          irqarray11_nc_b11s121;
wire          irqarray11_nc_b11s131;
wire          irqarray11_nc_b11s141;
wire          irqarray11_nc_b11s151;
reg    [15:0] irqarray11_pending_status;
wire          irqarray11_pending_we;
reg           irqarray11_pending_re;
reg    [15:0] irqarray11_pending_r;
wire          irqarray11_i2s_rx_dupe2;
wire          irqarray11_i2s_tx_dupe2;
wire          irqarray11_nc_b11s22;
wire          irqarray11_nc_b11s32;
wire          irqarray11_nc_b11s42;
wire          irqarray11_nc_b11s52;
wire          irqarray11_nc_b11s62;
wire          irqarray11_nc_b11s72;
wire          irqarray11_nc_b11s82;
wire          irqarray11_nc_b11s92;
wire          irqarray11_nc_b11s102;
wire          irqarray11_nc_b11s112;
wire          irqarray11_nc_b11s122;
wire          irqarray11_nc_b11s132;
wire          irqarray11_nc_b11s142;
wire          irqarray11_nc_b11s152;
reg    [15:0] irqarray11_enable_storage;
reg           irqarray11_enable_re;
wire          irqarray12_irq;
wire   [15:0] irqarray12_interrupts;
reg    [15:0] irqarray12_trigger;
reg    [15:0] irqarray12_soft_storage;
reg           irqarray12_soft_re;
wire   [15:0] irqarray12_use_edge;
reg    [15:0] irqarray12_edge_triggered_storage;
reg           irqarray12_edge_triggered_re;
wire   [15:0] irqarray12_rising;
reg    [15:0] irqarray12_polarity_storage;
reg           irqarray12_polarity_re;
wire          irqarray12_eventsourceflex192_status;
reg           irqarray12_eventsourceflex192_pending;
reg           irqarray12_eventsourceflex192_clear;
reg           irqarray12_eventsourceflex192_trigger_d;
reg           irqarray12_eventsourceflex192_trigger_filtered;
wire          irqarray12_eventsourceflex193_status;
reg           irqarray12_eventsourceflex193_pending;
reg           irqarray12_eventsourceflex193_clear;
reg           irqarray12_eventsourceflex193_trigger_d;
reg           irqarray12_eventsourceflex193_trigger_filtered;
wire          irqarray12_eventsourceflex194_status;
reg           irqarray12_eventsourceflex194_pending;
reg           irqarray12_eventsourceflex194_clear;
reg           irqarray12_eventsourceflex194_trigger_d;
reg           irqarray12_eventsourceflex194_trigger_filtered;
wire          irqarray12_eventsourceflex195_status;
reg           irqarray12_eventsourceflex195_pending;
reg           irqarray12_eventsourceflex195_clear;
reg           irqarray12_eventsourceflex195_trigger_d;
reg           irqarray12_eventsourceflex195_trigger_filtered;
wire          irqarray12_eventsourceflex196_status;
reg           irqarray12_eventsourceflex196_pending;
reg           irqarray12_eventsourceflex196_clear;
reg           irqarray12_eventsourceflex196_trigger_d;
reg           irqarray12_eventsourceflex196_trigger_filtered;
wire          irqarray12_eventsourceflex197_status;
reg           irqarray12_eventsourceflex197_pending;
reg           irqarray12_eventsourceflex197_clear;
reg           irqarray12_eventsourceflex197_trigger_d;
reg           irqarray12_eventsourceflex197_trigger_filtered;
wire          irqarray12_eventsourceflex198_status;
reg           irqarray12_eventsourceflex198_pending;
reg           irqarray12_eventsourceflex198_clear;
reg           irqarray12_eventsourceflex198_trigger_d;
reg           irqarray12_eventsourceflex198_trigger_filtered;
wire          irqarray12_eventsourceflex199_status;
reg           irqarray12_eventsourceflex199_pending;
reg           irqarray12_eventsourceflex199_clear;
reg           irqarray12_eventsourceflex199_trigger_d;
reg           irqarray12_eventsourceflex199_trigger_filtered;
wire          irqarray12_eventsourceflex200_status;
reg           irqarray12_eventsourceflex200_pending;
reg           irqarray12_eventsourceflex200_clear;
reg           irqarray12_eventsourceflex200_trigger_d;
reg           irqarray12_eventsourceflex200_trigger_filtered;
wire          irqarray12_eventsourceflex201_status;
reg           irqarray12_eventsourceflex201_pending;
reg           irqarray12_eventsourceflex201_clear;
reg           irqarray12_eventsourceflex201_trigger_d;
reg           irqarray12_eventsourceflex201_trigger_filtered;
wire          irqarray12_eventsourceflex202_status;
reg           irqarray12_eventsourceflex202_pending;
reg           irqarray12_eventsourceflex202_clear;
reg           irqarray12_eventsourceflex202_trigger_d;
reg           irqarray12_eventsourceflex202_trigger_filtered;
wire          irqarray12_eventsourceflex203_status;
reg           irqarray12_eventsourceflex203_pending;
reg           irqarray12_eventsourceflex203_clear;
reg           irqarray12_eventsourceflex203_trigger_d;
reg           irqarray12_eventsourceflex203_trigger_filtered;
wire          irqarray12_eventsourceflex204_status;
reg           irqarray12_eventsourceflex204_pending;
reg           irqarray12_eventsourceflex204_clear;
reg           irqarray12_eventsourceflex204_trigger_d;
reg           irqarray12_eventsourceflex204_trigger_filtered;
wire          irqarray12_eventsourceflex205_status;
reg           irqarray12_eventsourceflex205_pending;
reg           irqarray12_eventsourceflex205_clear;
reg           irqarray12_eventsourceflex205_trigger_d;
reg           irqarray12_eventsourceflex205_trigger_filtered;
wire          irqarray12_eventsourceflex206_status;
reg           irqarray12_eventsourceflex206_pending;
reg           irqarray12_eventsourceflex206_clear;
reg           irqarray12_eventsourceflex206_trigger_d;
reg           irqarray12_eventsourceflex206_trigger_filtered;
wire          irqarray12_eventsourceflex207_status;
reg           irqarray12_eventsourceflex207_pending;
reg           irqarray12_eventsourceflex207_clear;
reg           irqarray12_eventsourceflex207_trigger_d;
reg           irqarray12_eventsourceflex207_trigger_filtered;
wire          irqarray12_nc_b12s00;
wire          irqarray12_nc_b12s10;
wire          irqarray12_nc_b12s20;
wire          irqarray12_nc_b12s30;
wire          irqarray12_nc_b12s40;
wire          irqarray12_nc_b12s50;
wire          irqarray12_nc_b12s60;
wire          irqarray12_nc_b12s70;
wire          irqarray12_i2c0_nack0;
wire          irqarray12_i2c1_nack0;
wire          irqarray12_i2c2_nack0;
wire          irqarray12_i2c3_nack0;
wire          irqarray12_i2c0_err0;
wire          irqarray12_i2c1_err0;
wire          irqarray12_i2c2_err0;
wire          irqarray12_i2c3_err0;
reg    [15:0] irqarray12_status_status;
wire          irqarray12_status_we;
reg           irqarray12_status_re;
wire          irqarray12_nc_b12s01;
wire          irqarray12_nc_b12s11;
wire          irqarray12_nc_b12s21;
wire          irqarray12_nc_b12s31;
wire          irqarray12_nc_b12s41;
wire          irqarray12_nc_b12s51;
wire          irqarray12_nc_b12s61;
wire          irqarray12_nc_b12s71;
wire          irqarray12_i2c0_nack1;
wire          irqarray12_i2c1_nack1;
wire          irqarray12_i2c2_nack1;
wire          irqarray12_i2c3_nack1;
wire          irqarray12_i2c0_err1;
wire          irqarray12_i2c1_err1;
wire          irqarray12_i2c2_err1;
wire          irqarray12_i2c3_err1;
reg    [15:0] irqarray12_pending_status;
wire          irqarray12_pending_we;
reg           irqarray12_pending_re;
reg    [15:0] irqarray12_pending_r;
wire          irqarray12_nc_b12s02;
wire          irqarray12_nc_b12s12;
wire          irqarray12_nc_b12s22;
wire          irqarray12_nc_b12s32;
wire          irqarray12_nc_b12s42;
wire          irqarray12_nc_b12s52;
wire          irqarray12_nc_b12s62;
wire          irqarray12_nc_b12s72;
wire          irqarray12_i2c0_nack2;
wire          irqarray12_i2c1_nack2;
wire          irqarray12_i2c2_nack2;
wire          irqarray12_i2c3_nack2;
wire          irqarray12_i2c0_err2;
wire          irqarray12_i2c1_err2;
wire          irqarray12_i2c2_err2;
wire          irqarray12_i2c3_err2;
reg    [15:0] irqarray12_enable_storage;
reg           irqarray12_enable_re;
wire          irqarray13_irq;
wire   [15:0] irqarray13_interrupts;
reg    [15:0] irqarray13_trigger;
reg    [15:0] irqarray13_soft_storage;
reg           irqarray13_soft_re;
wire   [15:0] irqarray13_use_edge;
reg    [15:0] irqarray13_edge_triggered_storage;
reg           irqarray13_edge_triggered_re;
wire   [15:0] irqarray13_rising;
reg    [15:0] irqarray13_polarity_storage;
reg           irqarray13_polarity_re;
wire          irqarray13_eventsourceflex208_status;
reg           irqarray13_eventsourceflex208_pending;
reg           irqarray13_eventsourceflex208_clear;
reg           irqarray13_eventsourceflex208_trigger_d;
reg           irqarray13_eventsourceflex208_trigger_filtered;
wire          irqarray13_eventsourceflex209_status;
reg           irqarray13_eventsourceflex209_pending;
reg           irqarray13_eventsourceflex209_clear;
reg           irqarray13_eventsourceflex209_trigger_d;
reg           irqarray13_eventsourceflex209_trigger_filtered;
wire          irqarray13_eventsourceflex210_status;
reg           irqarray13_eventsourceflex210_pending;
reg           irqarray13_eventsourceflex210_clear;
reg           irqarray13_eventsourceflex210_trigger_d;
reg           irqarray13_eventsourceflex210_trigger_filtered;
wire          irqarray13_eventsourceflex211_status;
reg           irqarray13_eventsourceflex211_pending;
reg           irqarray13_eventsourceflex211_clear;
reg           irqarray13_eventsourceflex211_trigger_d;
reg           irqarray13_eventsourceflex211_trigger_filtered;
wire          irqarray13_eventsourceflex212_status;
reg           irqarray13_eventsourceflex212_pending;
reg           irqarray13_eventsourceflex212_clear;
reg           irqarray13_eventsourceflex212_trigger_d;
reg           irqarray13_eventsourceflex212_trigger_filtered;
wire          irqarray13_eventsourceflex213_status;
reg           irqarray13_eventsourceflex213_pending;
reg           irqarray13_eventsourceflex213_clear;
reg           irqarray13_eventsourceflex213_trigger_d;
reg           irqarray13_eventsourceflex213_trigger_filtered;
wire          irqarray13_eventsourceflex214_status;
reg           irqarray13_eventsourceflex214_pending;
reg           irqarray13_eventsourceflex214_clear;
reg           irqarray13_eventsourceflex214_trigger_d;
reg           irqarray13_eventsourceflex214_trigger_filtered;
wire          irqarray13_eventsourceflex215_status;
reg           irqarray13_eventsourceflex215_pending;
reg           irqarray13_eventsourceflex215_clear;
reg           irqarray13_eventsourceflex215_trigger_d;
reg           irqarray13_eventsourceflex215_trigger_filtered;
wire          irqarray13_eventsourceflex216_status;
reg           irqarray13_eventsourceflex216_pending;
reg           irqarray13_eventsourceflex216_clear;
reg           irqarray13_eventsourceflex216_trigger_d;
reg           irqarray13_eventsourceflex216_trigger_filtered;
wire          irqarray13_eventsourceflex217_status;
reg           irqarray13_eventsourceflex217_pending;
reg           irqarray13_eventsourceflex217_clear;
reg           irqarray13_eventsourceflex217_trigger_d;
reg           irqarray13_eventsourceflex217_trigger_filtered;
wire          irqarray13_eventsourceflex218_status;
reg           irqarray13_eventsourceflex218_pending;
reg           irqarray13_eventsourceflex218_clear;
reg           irqarray13_eventsourceflex218_trigger_d;
reg           irqarray13_eventsourceflex218_trigger_filtered;
wire          irqarray13_eventsourceflex219_status;
reg           irqarray13_eventsourceflex219_pending;
reg           irqarray13_eventsourceflex219_clear;
reg           irqarray13_eventsourceflex219_trigger_d;
reg           irqarray13_eventsourceflex219_trigger_filtered;
wire          irqarray13_eventsourceflex220_status;
reg           irqarray13_eventsourceflex220_pending;
reg           irqarray13_eventsourceflex220_clear;
reg           irqarray13_eventsourceflex220_trigger_d;
reg           irqarray13_eventsourceflex220_trigger_filtered;
wire          irqarray13_eventsourceflex221_status;
reg           irqarray13_eventsourceflex221_pending;
reg           irqarray13_eventsourceflex221_clear;
reg           irqarray13_eventsourceflex221_trigger_d;
reg           irqarray13_eventsourceflex221_trigger_filtered;
wire          irqarray13_eventsourceflex222_status;
reg           irqarray13_eventsourceflex222_pending;
reg           irqarray13_eventsourceflex222_clear;
reg           irqarray13_eventsourceflex222_trigger_d;
reg           irqarray13_eventsourceflex222_trigger_filtered;
wire          irqarray13_eventsourceflex223_status;
reg           irqarray13_eventsourceflex223_pending;
reg           irqarray13_eventsourceflex223_clear;
reg           irqarray13_eventsourceflex223_trigger_d;
reg           irqarray13_eventsourceflex223_trigger_filtered;
wire          irqarray13_coresuberr0;
wire          irqarray13_sceerr0;
wire          irqarray13_ifsuberr0;
wire          irqarray13_secirq0;
wire          irqarray13_nc_b13s40;
wire          irqarray13_nc_b13s50;
wire          irqarray13_nc_b13s60;
wire          irqarray13_nc_b13s70;
wire          irqarray13_nc_b13s80;
wire          irqarray13_nc_b13s90;
wire          irqarray13_nc_b13s100;
wire          irqarray13_nc_b13s110;
wire          irqarray13_nc_b13s120;
wire          irqarray13_nc_b13s130;
wire          irqarray13_nc_b13s140;
wire          irqarray13_nc_b13s150;
reg    [15:0] irqarray13_status_status;
wire          irqarray13_status_we;
reg           irqarray13_status_re;
wire          irqarray13_coresuberr1;
wire          irqarray13_sceerr1;
wire          irqarray13_ifsuberr1;
wire          irqarray13_secirq1;
wire          irqarray13_nc_b13s41;
wire          irqarray13_nc_b13s51;
wire          irqarray13_nc_b13s61;
wire          irqarray13_nc_b13s71;
wire          irqarray13_nc_b13s81;
wire          irqarray13_nc_b13s91;
wire          irqarray13_nc_b13s101;
wire          irqarray13_nc_b13s111;
wire          irqarray13_nc_b13s121;
wire          irqarray13_nc_b13s131;
wire          irqarray13_nc_b13s141;
wire          irqarray13_nc_b13s151;
reg    [15:0] irqarray13_pending_status;
wire          irqarray13_pending_we;
reg           irqarray13_pending_re;
reg    [15:0] irqarray13_pending_r;
wire          irqarray13_coresuberr2;
wire          irqarray13_sceerr2;
wire          irqarray13_ifsuberr2;
wire          irqarray13_secirq2;
wire          irqarray13_nc_b13s42;
wire          irqarray13_nc_b13s52;
wire          irqarray13_nc_b13s62;
wire          irqarray13_nc_b13s72;
wire          irqarray13_nc_b13s82;
wire          irqarray13_nc_b13s92;
wire          irqarray13_nc_b13s102;
wire          irqarray13_nc_b13s112;
wire          irqarray13_nc_b13s122;
wire          irqarray13_nc_b13s132;
wire          irqarray13_nc_b13s142;
wire          irqarray13_nc_b13s152;
reg    [15:0] irqarray13_enable_storage;
reg           irqarray13_enable_re;
wire          irqarray14_irq;
wire   [15:0] irqarray14_interrupts;
reg    [15:0] irqarray14_trigger;
reg    [15:0] irqarray14_soft_storage;
reg           irqarray14_soft_re;
wire   [15:0] irqarray14_use_edge;
reg    [15:0] irqarray14_edge_triggered_storage;
reg           irqarray14_edge_triggered_re;
wire   [15:0] irqarray14_rising;
reg    [15:0] irqarray14_polarity_storage;
reg           irqarray14_polarity_re;
wire          irqarray14_eventsourceflex224_status;
reg           irqarray14_eventsourceflex224_pending;
reg           irqarray14_eventsourceflex224_clear;
reg           irqarray14_eventsourceflex224_trigger_d;
reg           irqarray14_eventsourceflex224_trigger_filtered;
wire          irqarray14_eventsourceflex225_status;
reg           irqarray14_eventsourceflex225_pending;
reg           irqarray14_eventsourceflex225_clear;
reg           irqarray14_eventsourceflex225_trigger_d;
reg           irqarray14_eventsourceflex225_trigger_filtered;
wire          irqarray14_eventsourceflex226_status;
reg           irqarray14_eventsourceflex226_pending;
reg           irqarray14_eventsourceflex226_clear;
reg           irqarray14_eventsourceflex226_trigger_d;
reg           irqarray14_eventsourceflex226_trigger_filtered;
wire          irqarray14_eventsourceflex227_status;
reg           irqarray14_eventsourceflex227_pending;
reg           irqarray14_eventsourceflex227_clear;
reg           irqarray14_eventsourceflex227_trigger_d;
reg           irqarray14_eventsourceflex227_trigger_filtered;
wire          irqarray14_eventsourceflex228_status;
reg           irqarray14_eventsourceflex228_pending;
reg           irqarray14_eventsourceflex228_clear;
reg           irqarray14_eventsourceflex228_trigger_d;
reg           irqarray14_eventsourceflex228_trigger_filtered;
wire          irqarray14_eventsourceflex229_status;
reg           irqarray14_eventsourceflex229_pending;
reg           irqarray14_eventsourceflex229_clear;
reg           irqarray14_eventsourceflex229_trigger_d;
reg           irqarray14_eventsourceflex229_trigger_filtered;
wire          irqarray14_eventsourceflex230_status;
reg           irqarray14_eventsourceflex230_pending;
reg           irqarray14_eventsourceflex230_clear;
reg           irqarray14_eventsourceflex230_trigger_d;
reg           irqarray14_eventsourceflex230_trigger_filtered;
wire          irqarray14_eventsourceflex231_status;
reg           irqarray14_eventsourceflex231_pending;
reg           irqarray14_eventsourceflex231_clear;
reg           irqarray14_eventsourceflex231_trigger_d;
reg           irqarray14_eventsourceflex231_trigger_filtered;
wire          irqarray14_eventsourceflex232_status;
reg           irqarray14_eventsourceflex232_pending;
reg           irqarray14_eventsourceflex232_clear;
reg           irqarray14_eventsourceflex232_trigger_d;
reg           irqarray14_eventsourceflex232_trigger_filtered;
wire          irqarray14_eventsourceflex233_status;
reg           irqarray14_eventsourceflex233_pending;
reg           irqarray14_eventsourceflex233_clear;
reg           irqarray14_eventsourceflex233_trigger_d;
reg           irqarray14_eventsourceflex233_trigger_filtered;
wire          irqarray14_eventsourceflex234_status;
reg           irqarray14_eventsourceflex234_pending;
reg           irqarray14_eventsourceflex234_clear;
reg           irqarray14_eventsourceflex234_trigger_d;
reg           irqarray14_eventsourceflex234_trigger_filtered;
wire          irqarray14_eventsourceflex235_status;
reg           irqarray14_eventsourceflex235_pending;
reg           irqarray14_eventsourceflex235_clear;
reg           irqarray14_eventsourceflex235_trigger_d;
reg           irqarray14_eventsourceflex235_trigger_filtered;
wire          irqarray14_eventsourceflex236_status;
reg           irqarray14_eventsourceflex236_pending;
reg           irqarray14_eventsourceflex236_clear;
reg           irqarray14_eventsourceflex236_trigger_d;
reg           irqarray14_eventsourceflex236_trigger_filtered;
wire          irqarray14_eventsourceflex237_status;
reg           irqarray14_eventsourceflex237_pending;
reg           irqarray14_eventsourceflex237_clear;
reg           irqarray14_eventsourceflex237_trigger_d;
reg           irqarray14_eventsourceflex237_trigger_filtered;
wire          irqarray14_eventsourceflex238_status;
reg           irqarray14_eventsourceflex238_pending;
reg           irqarray14_eventsourceflex238_clear;
reg           irqarray14_eventsourceflex238_trigger_d;
reg           irqarray14_eventsourceflex238_trigger_filtered;
wire          irqarray14_eventsourceflex239_status;
reg           irqarray14_eventsourceflex239_pending;
reg           irqarray14_eventsourceflex239_clear;
reg           irqarray14_eventsourceflex239_trigger_d;
reg           irqarray14_eventsourceflex239_trigger_filtered;
wire          irqarray14_uart2_rx_dupe0;
wire          irqarray14_uart2_tx_dupe0;
wire          irqarray14_uart2_rx_char_dupe0;
wire          irqarray14_uart2_err_dupe0;
wire          irqarray14_uart3_rx_dupe0;
wire          irqarray14_uart3_tx_dupe0;
wire          irqarray14_uart3_rx_char_dupe0;
wire          irqarray14_uart3_err_dupe0;
wire          irqarray14_trng_done_dupe0;
wire          irqarray14_nc_b14s90;
wire          irqarray14_nc_b14s100;
wire          irqarray14_nc_b14s110;
wire          irqarray14_nc_b14s120;
wire          irqarray14_nc_b14s130;
wire          irqarray14_nc_b14s140;
wire          irqarray14_nc_b14s150;
reg    [15:0] irqarray14_status_status;
wire          irqarray14_status_we;
reg           irqarray14_status_re;
wire          irqarray14_uart2_rx_dupe1;
wire          irqarray14_uart2_tx_dupe1;
wire          irqarray14_uart2_rx_char_dupe1;
wire          irqarray14_uart2_err_dupe1;
wire          irqarray14_uart3_rx_dupe1;
wire          irqarray14_uart3_tx_dupe1;
wire          irqarray14_uart3_rx_char_dupe1;
wire          irqarray14_uart3_err_dupe1;
wire          irqarray14_trng_done_dupe1;
wire          irqarray14_nc_b14s91;
wire          irqarray14_nc_b14s101;
wire          irqarray14_nc_b14s111;
wire          irqarray14_nc_b14s121;
wire          irqarray14_nc_b14s131;
wire          irqarray14_nc_b14s141;
wire          irqarray14_nc_b14s151;
reg    [15:0] irqarray14_pending_status;
wire          irqarray14_pending_we;
reg           irqarray14_pending_re;
reg    [15:0] irqarray14_pending_r;
wire          irqarray14_uart2_rx_dupe2;
wire          irqarray14_uart2_tx_dupe2;
wire          irqarray14_uart2_rx_char_dupe2;
wire          irqarray14_uart2_err_dupe2;
wire          irqarray14_uart3_rx_dupe2;
wire          irqarray14_uart3_tx_dupe2;
wire          irqarray14_uart3_rx_char_dupe2;
wire          irqarray14_uart3_err_dupe2;
wire          irqarray14_trng_done_dupe2;
wire          irqarray14_nc_b14s92;
wire          irqarray14_nc_b14s102;
wire          irqarray14_nc_b14s112;
wire          irqarray14_nc_b14s122;
wire          irqarray14_nc_b14s132;
wire          irqarray14_nc_b14s142;
wire          irqarray14_nc_b14s152;
reg    [15:0] irqarray14_enable_storage;
reg           irqarray14_enable_re;
wire          irqarray15_irq;
wire   [15:0] irqarray15_interrupts;
reg    [15:0] irqarray15_trigger;
reg    [15:0] irqarray15_soft_storage;
reg           irqarray15_soft_re;
wire   [15:0] irqarray15_use_edge;
reg    [15:0] irqarray15_edge_triggered_storage;
reg           irqarray15_edge_triggered_re;
wire   [15:0] irqarray15_rising;
reg    [15:0] irqarray15_polarity_storage;
reg           irqarray15_polarity_re;
wire          irqarray15_eventsourceflex240_status;
reg           irqarray15_eventsourceflex240_pending;
reg           irqarray15_eventsourceflex240_clear;
reg           irqarray15_eventsourceflex240_trigger_d;
reg           irqarray15_eventsourceflex240_trigger_filtered;
wire          irqarray15_eventsourceflex241_status;
reg           irqarray15_eventsourceflex241_pending;
reg           irqarray15_eventsourceflex241_clear;
reg           irqarray15_eventsourceflex241_trigger_d;
reg           irqarray15_eventsourceflex241_trigger_filtered;
wire          irqarray15_eventsourceflex242_status;
reg           irqarray15_eventsourceflex242_pending;
reg           irqarray15_eventsourceflex242_clear;
reg           irqarray15_eventsourceflex242_trigger_d;
reg           irqarray15_eventsourceflex242_trigger_filtered;
wire          irqarray15_eventsourceflex243_status;
reg           irqarray15_eventsourceflex243_pending;
reg           irqarray15_eventsourceflex243_clear;
reg           irqarray15_eventsourceflex243_trigger_d;
reg           irqarray15_eventsourceflex243_trigger_filtered;
wire          irqarray15_eventsourceflex244_status;
reg           irqarray15_eventsourceflex244_pending;
reg           irqarray15_eventsourceflex244_clear;
reg           irqarray15_eventsourceflex244_trigger_d;
reg           irqarray15_eventsourceflex244_trigger_filtered;
wire          irqarray15_eventsourceflex245_status;
reg           irqarray15_eventsourceflex245_pending;
reg           irqarray15_eventsourceflex245_clear;
reg           irqarray15_eventsourceflex245_trigger_d;
reg           irqarray15_eventsourceflex245_trigger_filtered;
wire          irqarray15_eventsourceflex246_status;
reg           irqarray15_eventsourceflex246_pending;
reg           irqarray15_eventsourceflex246_clear;
reg           irqarray15_eventsourceflex246_trigger_d;
reg           irqarray15_eventsourceflex246_trigger_filtered;
wire          irqarray15_eventsourceflex247_status;
reg           irqarray15_eventsourceflex247_pending;
reg           irqarray15_eventsourceflex247_clear;
reg           irqarray15_eventsourceflex247_trigger_d;
reg           irqarray15_eventsourceflex247_trigger_filtered;
wire          irqarray15_eventsourceflex248_status;
reg           irqarray15_eventsourceflex248_pending;
reg           irqarray15_eventsourceflex248_clear;
reg           irqarray15_eventsourceflex248_trigger_d;
reg           irqarray15_eventsourceflex248_trigger_filtered;
wire          irqarray15_eventsourceflex249_status;
reg           irqarray15_eventsourceflex249_pending;
reg           irqarray15_eventsourceflex249_clear;
reg           irqarray15_eventsourceflex249_trigger_d;
reg           irqarray15_eventsourceflex249_trigger_filtered;
wire          irqarray15_eventsourceflex250_status;
reg           irqarray15_eventsourceflex250_pending;
reg           irqarray15_eventsourceflex250_clear;
reg           irqarray15_eventsourceflex250_trigger_d;
reg           irqarray15_eventsourceflex250_trigger_filtered;
wire          irqarray15_eventsourceflex251_status;
reg           irqarray15_eventsourceflex251_pending;
reg           irqarray15_eventsourceflex251_clear;
reg           irqarray15_eventsourceflex251_trigger_d;
reg           irqarray15_eventsourceflex251_trigger_filtered;
wire          irqarray15_eventsourceflex252_status;
reg           irqarray15_eventsourceflex252_pending;
reg           irqarray15_eventsourceflex252_clear;
reg           irqarray15_eventsourceflex252_trigger_d;
reg           irqarray15_eventsourceflex252_trigger_filtered;
wire          irqarray15_eventsourceflex253_status;
reg           irqarray15_eventsourceflex253_pending;
reg           irqarray15_eventsourceflex253_clear;
reg           irqarray15_eventsourceflex253_trigger_d;
reg           irqarray15_eventsourceflex253_trigger_filtered;
wire          irqarray15_eventsourceflex254_status;
reg           irqarray15_eventsourceflex254_pending;
reg           irqarray15_eventsourceflex254_clear;
reg           irqarray15_eventsourceflex254_trigger_d;
reg           irqarray15_eventsourceflex254_trigger_filtered;
wire          irqarray15_eventsourceflex255_status;
reg           irqarray15_eventsourceflex255_pending;
reg           irqarray15_eventsourceflex255_clear;
reg           irqarray15_eventsourceflex255_trigger_d;
reg           irqarray15_eventsourceflex255_trigger_filtered;
wire          irqarray15_sec00;
wire          irqarray15_nc_b15s10;
wire          irqarray15_nc_b15s20;
wire          irqarray15_nc_b15s30;
wire          irqarray15_nc_b15s40;
wire          irqarray15_nc_b15s50;
wire          irqarray15_nc_b15s60;
wire          irqarray15_nc_b15s70;
wire          irqarray15_nc_b15s80;
wire          irqarray15_nc_b15s90;
wire          irqarray15_nc_b15s100;
wire          irqarray15_nc_b15s110;
wire          irqarray15_nc_b15s120;
wire          irqarray15_nc_b15s130;
wire          irqarray15_nc_b15s140;
wire          irqarray15_nc_b15s150;
reg    [15:0] irqarray15_status_status;
wire          irqarray15_status_we;
reg           irqarray15_status_re;
wire          irqarray15_sec01;
wire          irqarray15_nc_b15s11;
wire          irqarray15_nc_b15s21;
wire          irqarray15_nc_b15s31;
wire          irqarray15_nc_b15s41;
wire          irqarray15_nc_b15s51;
wire          irqarray15_nc_b15s61;
wire          irqarray15_nc_b15s71;
wire          irqarray15_nc_b15s81;
wire          irqarray15_nc_b15s91;
wire          irqarray15_nc_b15s101;
wire          irqarray15_nc_b15s111;
wire          irqarray15_nc_b15s121;
wire          irqarray15_nc_b15s131;
wire          irqarray15_nc_b15s141;
wire          irqarray15_nc_b15s151;
reg    [15:0] irqarray15_pending_status;
wire          irqarray15_pending_we;
reg           irqarray15_pending_re;
reg    [15:0] irqarray15_pending_r;
wire          irqarray15_sec02;
wire          irqarray15_nc_b15s12;
wire          irqarray15_nc_b15s22;
wire          irqarray15_nc_b15s32;
wire          irqarray15_nc_b15s42;
wire          irqarray15_nc_b15s52;
wire          irqarray15_nc_b15s62;
wire          irqarray15_nc_b15s72;
wire          irqarray15_nc_b15s82;
wire          irqarray15_nc_b15s92;
wire          irqarray15_nc_b15s102;
wire          irqarray15_nc_b15s112;
wire          irqarray15_nc_b15s122;
wire          irqarray15_nc_b15s132;
wire          irqarray15_nc_b15s142;
wire          irqarray15_nc_b15s152;
reg    [15:0] irqarray15_enable_storage;
reg           irqarray15_enable_re;
wire          irqarray16_irq;
wire   [15:0] irqarray16_interrupts;
reg    [15:0] irqarray16_trigger;
reg    [15:0] irqarray16_soft_storage;
reg           irqarray16_soft_re;
wire   [15:0] irqarray16_use_edge;
reg    [15:0] irqarray16_edge_triggered_storage;
reg           irqarray16_edge_triggered_re;
wire   [15:0] irqarray16_rising;
reg    [15:0] irqarray16_polarity_storage;
reg           irqarray16_polarity_re;
wire          irqarray16_eventsourceflex256_status;
reg           irqarray16_eventsourceflex256_pending;
reg           irqarray16_eventsourceflex256_clear;
reg           irqarray16_eventsourceflex256_trigger_d;
reg           irqarray16_eventsourceflex256_trigger_filtered;
wire          irqarray16_eventsourceflex257_status;
reg           irqarray16_eventsourceflex257_pending;
reg           irqarray16_eventsourceflex257_clear;
reg           irqarray16_eventsourceflex257_trigger_d;
reg           irqarray16_eventsourceflex257_trigger_filtered;
wire          irqarray16_eventsourceflex258_status;
reg           irqarray16_eventsourceflex258_pending;
reg           irqarray16_eventsourceflex258_clear;
reg           irqarray16_eventsourceflex258_trigger_d;
reg           irqarray16_eventsourceflex258_trigger_filtered;
wire          irqarray16_eventsourceflex259_status;
reg           irqarray16_eventsourceflex259_pending;
reg           irqarray16_eventsourceflex259_clear;
reg           irqarray16_eventsourceflex259_trigger_d;
reg           irqarray16_eventsourceflex259_trigger_filtered;
wire          irqarray16_eventsourceflex260_status;
reg           irqarray16_eventsourceflex260_pending;
reg           irqarray16_eventsourceflex260_clear;
reg           irqarray16_eventsourceflex260_trigger_d;
reg           irqarray16_eventsourceflex260_trigger_filtered;
wire          irqarray16_eventsourceflex261_status;
reg           irqarray16_eventsourceflex261_pending;
reg           irqarray16_eventsourceflex261_clear;
reg           irqarray16_eventsourceflex261_trigger_d;
reg           irqarray16_eventsourceflex261_trigger_filtered;
wire          irqarray16_eventsourceflex262_status;
reg           irqarray16_eventsourceflex262_pending;
reg           irqarray16_eventsourceflex262_clear;
reg           irqarray16_eventsourceflex262_trigger_d;
reg           irqarray16_eventsourceflex262_trigger_filtered;
wire          irqarray16_eventsourceflex263_status;
reg           irqarray16_eventsourceflex263_pending;
reg           irqarray16_eventsourceflex263_clear;
reg           irqarray16_eventsourceflex263_trigger_d;
reg           irqarray16_eventsourceflex263_trigger_filtered;
wire          irqarray16_eventsourceflex264_status;
reg           irqarray16_eventsourceflex264_pending;
reg           irqarray16_eventsourceflex264_clear;
reg           irqarray16_eventsourceflex264_trigger_d;
reg           irqarray16_eventsourceflex264_trigger_filtered;
wire          irqarray16_eventsourceflex265_status;
reg           irqarray16_eventsourceflex265_pending;
reg           irqarray16_eventsourceflex265_clear;
reg           irqarray16_eventsourceflex265_trigger_d;
reg           irqarray16_eventsourceflex265_trigger_filtered;
wire          irqarray16_eventsourceflex266_status;
reg           irqarray16_eventsourceflex266_pending;
reg           irqarray16_eventsourceflex266_clear;
reg           irqarray16_eventsourceflex266_trigger_d;
reg           irqarray16_eventsourceflex266_trigger_filtered;
wire          irqarray16_eventsourceflex267_status;
reg           irqarray16_eventsourceflex267_pending;
reg           irqarray16_eventsourceflex267_clear;
reg           irqarray16_eventsourceflex267_trigger_d;
reg           irqarray16_eventsourceflex267_trigger_filtered;
wire          irqarray16_eventsourceflex268_status;
reg           irqarray16_eventsourceflex268_pending;
reg           irqarray16_eventsourceflex268_clear;
reg           irqarray16_eventsourceflex268_trigger_d;
reg           irqarray16_eventsourceflex268_trigger_filtered;
wire          irqarray16_eventsourceflex269_status;
reg           irqarray16_eventsourceflex269_pending;
reg           irqarray16_eventsourceflex269_clear;
reg           irqarray16_eventsourceflex269_trigger_d;
reg           irqarray16_eventsourceflex269_trigger_filtered;
wire          irqarray16_eventsourceflex270_status;
reg           irqarray16_eventsourceflex270_pending;
reg           irqarray16_eventsourceflex270_clear;
reg           irqarray16_eventsourceflex270_trigger_d;
reg           irqarray16_eventsourceflex270_trigger_filtered;
wire          irqarray16_eventsourceflex271_status;
reg           irqarray16_eventsourceflex271_pending;
reg           irqarray16_eventsourceflex271_clear;
reg           irqarray16_eventsourceflex271_trigger_d;
reg           irqarray16_eventsourceflex271_trigger_filtered;
wire          irqarray16_cam_rx_dupe0;
wire          irqarray16_i2s_rx_dupe0;
wire          irqarray16_i2s_tx_dupe0;
wire          irqarray16_nc_b16s30;
wire          irqarray16_spim1_rx_dupe0;
wire          irqarray16_spim1_tx_dupe0;
wire          irqarray16_spim1_cmd_dupe0;
wire          irqarray16_spim1_eot_dupe0;
wire          irqarray16_spim2_rx_dupe0;
wire          irqarray16_spim2_tx_dupe0;
wire          irqarray16_spim2_cmd_dupe0;
wire          irqarray16_spim2_eot_dupe0;
wire          irqarray16_i2c0_rx_dupe0;
wire          irqarray16_i2c0_tx_dupe0;
wire          irqarray16_i2c0_cmd_dupe0;
wire          irqarray16_i2c0_eot_dupe0;
reg    [15:0] irqarray16_status_status;
wire          irqarray16_status_we;
reg           irqarray16_status_re;
wire          irqarray16_cam_rx_dupe1;
wire          irqarray16_i2s_rx_dupe1;
wire          irqarray16_i2s_tx_dupe1;
wire          irqarray16_nc_b16s31;
wire          irqarray16_spim1_rx_dupe1;
wire          irqarray16_spim1_tx_dupe1;
wire          irqarray16_spim1_cmd_dupe1;
wire          irqarray16_spim1_eot_dupe1;
wire          irqarray16_spim2_rx_dupe1;
wire          irqarray16_spim2_tx_dupe1;
wire          irqarray16_spim2_cmd_dupe1;
wire          irqarray16_spim2_eot_dupe1;
wire          irqarray16_i2c0_rx_dupe1;
wire          irqarray16_i2c0_tx_dupe1;
wire          irqarray16_i2c0_cmd_dupe1;
wire          irqarray16_i2c0_eot_dupe1;
reg    [15:0] irqarray16_pending_status;
wire          irqarray16_pending_we;
reg           irqarray16_pending_re;
reg    [15:0] irqarray16_pending_r;
wire          irqarray16_cam_rx_dupe2;
wire          irqarray16_i2s_rx_dupe2;
wire          irqarray16_i2s_tx_dupe2;
wire          irqarray16_nc_b16s32;
wire          irqarray16_spim1_rx_dupe2;
wire          irqarray16_spim1_tx_dupe2;
wire          irqarray16_spim1_cmd_dupe2;
wire          irqarray16_spim1_eot_dupe2;
wire          irqarray16_spim2_rx_dupe2;
wire          irqarray16_spim2_tx_dupe2;
wire          irqarray16_spim2_cmd_dupe2;
wire          irqarray16_spim2_eot_dupe2;
wire          irqarray16_i2c0_rx_dupe2;
wire          irqarray16_i2c0_tx_dupe2;
wire          irqarray16_i2c0_cmd_dupe2;
wire          irqarray16_i2c0_eot_dupe2;
reg    [15:0] irqarray16_enable_storage;
reg           irqarray16_enable_re;
wire          irqarray17_irq;
wire   [15:0] irqarray17_interrupts;
reg    [15:0] irqarray17_trigger;
reg    [15:0] irqarray17_soft_storage;
reg           irqarray17_soft_re;
wire   [15:0] irqarray17_use_edge;
reg    [15:0] irqarray17_edge_triggered_storage;
reg           irqarray17_edge_triggered_re;
wire   [15:0] irqarray17_rising;
reg    [15:0] irqarray17_polarity_storage;
reg           irqarray17_polarity_re;
wire          irqarray17_eventsourceflex272_status;
reg           irqarray17_eventsourceflex272_pending;
reg           irqarray17_eventsourceflex272_clear;
reg           irqarray17_eventsourceflex272_trigger_d;
reg           irqarray17_eventsourceflex272_trigger_filtered;
wire          irqarray17_eventsourceflex273_status;
reg           irqarray17_eventsourceflex273_pending;
reg           irqarray17_eventsourceflex273_clear;
reg           irqarray17_eventsourceflex273_trigger_d;
reg           irqarray17_eventsourceflex273_trigger_filtered;
wire          irqarray17_eventsourceflex274_status;
reg           irqarray17_eventsourceflex274_pending;
reg           irqarray17_eventsourceflex274_clear;
reg           irqarray17_eventsourceflex274_trigger_d;
reg           irqarray17_eventsourceflex274_trigger_filtered;
wire          irqarray17_eventsourceflex275_status;
reg           irqarray17_eventsourceflex275_pending;
reg           irqarray17_eventsourceflex275_clear;
reg           irqarray17_eventsourceflex275_trigger_d;
reg           irqarray17_eventsourceflex275_trigger_filtered;
wire          irqarray17_eventsourceflex276_status;
reg           irqarray17_eventsourceflex276_pending;
reg           irqarray17_eventsourceflex276_clear;
reg           irqarray17_eventsourceflex276_trigger_d;
reg           irqarray17_eventsourceflex276_trigger_filtered;
wire          irqarray17_eventsourceflex277_status;
reg           irqarray17_eventsourceflex277_pending;
reg           irqarray17_eventsourceflex277_clear;
reg           irqarray17_eventsourceflex277_trigger_d;
reg           irqarray17_eventsourceflex277_trigger_filtered;
wire          irqarray17_eventsourceflex278_status;
reg           irqarray17_eventsourceflex278_pending;
reg           irqarray17_eventsourceflex278_clear;
reg           irqarray17_eventsourceflex278_trigger_d;
reg           irqarray17_eventsourceflex278_trigger_filtered;
wire          irqarray17_eventsourceflex279_status;
reg           irqarray17_eventsourceflex279_pending;
reg           irqarray17_eventsourceflex279_clear;
reg           irqarray17_eventsourceflex279_trigger_d;
reg           irqarray17_eventsourceflex279_trigger_filtered;
wire          irqarray17_eventsourceflex280_status;
reg           irqarray17_eventsourceflex280_pending;
reg           irqarray17_eventsourceflex280_clear;
reg           irqarray17_eventsourceflex280_trigger_d;
reg           irqarray17_eventsourceflex280_trigger_filtered;
wire          irqarray17_eventsourceflex281_status;
reg           irqarray17_eventsourceflex281_pending;
reg           irqarray17_eventsourceflex281_clear;
reg           irqarray17_eventsourceflex281_trigger_d;
reg           irqarray17_eventsourceflex281_trigger_filtered;
wire          irqarray17_eventsourceflex282_status;
reg           irqarray17_eventsourceflex282_pending;
reg           irqarray17_eventsourceflex282_clear;
reg           irqarray17_eventsourceflex282_trigger_d;
reg           irqarray17_eventsourceflex282_trigger_filtered;
wire          irqarray17_eventsourceflex283_status;
reg           irqarray17_eventsourceflex283_pending;
reg           irqarray17_eventsourceflex283_clear;
reg           irqarray17_eventsourceflex283_trigger_d;
reg           irqarray17_eventsourceflex283_trigger_filtered;
wire          irqarray17_eventsourceflex284_status;
reg           irqarray17_eventsourceflex284_pending;
reg           irqarray17_eventsourceflex284_clear;
reg           irqarray17_eventsourceflex284_trigger_d;
reg           irqarray17_eventsourceflex284_trigger_filtered;
wire          irqarray17_eventsourceflex285_status;
reg           irqarray17_eventsourceflex285_pending;
reg           irqarray17_eventsourceflex285_clear;
reg           irqarray17_eventsourceflex285_trigger_d;
reg           irqarray17_eventsourceflex285_trigger_filtered;
wire          irqarray17_eventsourceflex286_status;
reg           irqarray17_eventsourceflex286_pending;
reg           irqarray17_eventsourceflex286_clear;
reg           irqarray17_eventsourceflex286_trigger_d;
reg           irqarray17_eventsourceflex286_trigger_filtered;
wire          irqarray17_eventsourceflex287_status;
reg           irqarray17_eventsourceflex287_pending;
reg           irqarray17_eventsourceflex287_clear;
reg           irqarray17_eventsourceflex287_trigger_d;
reg           irqarray17_eventsourceflex287_trigger_filtered;
wire          irqarray17_i2c1_rx_dupe0;
wire          irqarray17_i2c1_tx_dupe0;
wire          irqarray17_i2c1_cmd_dupe0;
wire          irqarray17_i2c1_eot_dupe0;
wire          irqarray17_pioirq0_dupe0;
wire          irqarray17_pioirq1_dupe0;
wire          irqarray17_pioirq2_dupe0;
wire          irqarray17_pioirq3_dupe0;
wire          irqarray17_qfcirq_dupe0;
wire          irqarray17_adc_rx_dupe0;
wire          irqarray17_ioxirq_dupe0;
wire          irqarray17_sddcirq_dupe0;
wire          irqarray17_nc_b17s120;
wire          irqarray17_nc_b17s130;
wire          irqarray17_nc_b17s140;
wire          irqarray17_nc_b17s150;
reg    [15:0] irqarray17_status_status;
wire          irqarray17_status_we;
reg           irqarray17_status_re;
wire          irqarray17_i2c1_rx_dupe1;
wire          irqarray17_i2c1_tx_dupe1;
wire          irqarray17_i2c1_cmd_dupe1;
wire          irqarray17_i2c1_eot_dupe1;
wire          irqarray17_pioirq0_dupe1;
wire          irqarray17_pioirq1_dupe1;
wire          irqarray17_pioirq2_dupe1;
wire          irqarray17_pioirq3_dupe1;
wire          irqarray17_qfcirq_dupe1;
wire          irqarray17_adc_rx_dupe1;
wire          irqarray17_ioxirq_dupe1;
wire          irqarray17_sddcirq_dupe1;
wire          irqarray17_nc_b17s121;
wire          irqarray17_nc_b17s131;
wire          irqarray17_nc_b17s141;
wire          irqarray17_nc_b17s151;
reg    [15:0] irqarray17_pending_status;
wire          irqarray17_pending_we;
reg           irqarray17_pending_re;
reg    [15:0] irqarray17_pending_r;
wire          irqarray17_i2c1_rx_dupe2;
wire          irqarray17_i2c1_tx_dupe2;
wire          irqarray17_i2c1_cmd_dupe2;
wire          irqarray17_i2c1_eot_dupe2;
wire          irqarray17_pioirq0_dupe2;
wire          irqarray17_pioirq1_dupe2;
wire          irqarray17_pioirq2_dupe2;
wire          irqarray17_pioirq3_dupe2;
wire          irqarray17_qfcirq_dupe2;
wire          irqarray17_adc_rx_dupe2;
wire          irqarray17_ioxirq_dupe2;
wire          irqarray17_sddcirq_dupe2;
wire          irqarray17_nc_b17s122;
wire          irqarray17_nc_b17s132;
wire          irqarray17_nc_b17s142;
wire          irqarray17_nc_b17s152;
reg    [15:0] irqarray17_enable_storage;
reg           irqarray17_enable_re;
wire          irqarray18_irq;
wire   [15:0] irqarray18_interrupts;
reg    [15:0] irqarray18_trigger;
reg    [15:0] irqarray18_soft_storage;
reg           irqarray18_soft_re;
wire   [15:0] irqarray18_use_edge;
reg    [15:0] irqarray18_edge_triggered_storage;
reg           irqarray18_edge_triggered_re;
wire   [15:0] irqarray18_rising;
reg    [15:0] irqarray18_polarity_storage;
reg           irqarray18_polarity_re;
wire          irqarray18_eventsourceflex288_status;
reg           irqarray18_eventsourceflex288_pending;
reg           irqarray18_eventsourceflex288_clear;
reg           irqarray18_eventsourceflex288_trigger_d;
reg           irqarray18_eventsourceflex288_trigger_filtered;
wire          irqarray18_eventsourceflex289_status;
reg           irqarray18_eventsourceflex289_pending;
reg           irqarray18_eventsourceflex289_clear;
reg           irqarray18_eventsourceflex289_trigger_d;
reg           irqarray18_eventsourceflex289_trigger_filtered;
wire          irqarray18_eventsourceflex290_status;
reg           irqarray18_eventsourceflex290_pending;
reg           irqarray18_eventsourceflex290_clear;
reg           irqarray18_eventsourceflex290_trigger_d;
reg           irqarray18_eventsourceflex290_trigger_filtered;
wire          irqarray18_eventsourceflex291_status;
reg           irqarray18_eventsourceflex291_pending;
reg           irqarray18_eventsourceflex291_clear;
reg           irqarray18_eventsourceflex291_trigger_d;
reg           irqarray18_eventsourceflex291_trigger_filtered;
wire          irqarray18_eventsourceflex292_status;
reg           irqarray18_eventsourceflex292_pending;
reg           irqarray18_eventsourceflex292_clear;
reg           irqarray18_eventsourceflex292_trigger_d;
reg           irqarray18_eventsourceflex292_trigger_filtered;
wire          irqarray18_eventsourceflex293_status;
reg           irqarray18_eventsourceflex293_pending;
reg           irqarray18_eventsourceflex293_clear;
reg           irqarray18_eventsourceflex293_trigger_d;
reg           irqarray18_eventsourceflex293_trigger_filtered;
wire          irqarray18_eventsourceflex294_status;
reg           irqarray18_eventsourceflex294_pending;
reg           irqarray18_eventsourceflex294_clear;
reg           irqarray18_eventsourceflex294_trigger_d;
reg           irqarray18_eventsourceflex294_trigger_filtered;
wire          irqarray18_eventsourceflex295_status;
reg           irqarray18_eventsourceflex295_pending;
reg           irqarray18_eventsourceflex295_clear;
reg           irqarray18_eventsourceflex295_trigger_d;
reg           irqarray18_eventsourceflex295_trigger_filtered;
wire          irqarray18_eventsourceflex296_status;
reg           irqarray18_eventsourceflex296_pending;
reg           irqarray18_eventsourceflex296_clear;
reg           irqarray18_eventsourceflex296_trigger_d;
reg           irqarray18_eventsourceflex296_trigger_filtered;
wire          irqarray18_eventsourceflex297_status;
reg           irqarray18_eventsourceflex297_pending;
reg           irqarray18_eventsourceflex297_clear;
reg           irqarray18_eventsourceflex297_trigger_d;
reg           irqarray18_eventsourceflex297_trigger_filtered;
wire          irqarray18_eventsourceflex298_status;
reg           irqarray18_eventsourceflex298_pending;
reg           irqarray18_eventsourceflex298_clear;
reg           irqarray18_eventsourceflex298_trigger_d;
reg           irqarray18_eventsourceflex298_trigger_filtered;
wire          irqarray18_eventsourceflex299_status;
reg           irqarray18_eventsourceflex299_pending;
reg           irqarray18_eventsourceflex299_clear;
reg           irqarray18_eventsourceflex299_trigger_d;
reg           irqarray18_eventsourceflex299_trigger_filtered;
wire          irqarray18_eventsourceflex300_status;
reg           irqarray18_eventsourceflex300_pending;
reg           irqarray18_eventsourceflex300_clear;
reg           irqarray18_eventsourceflex300_trigger_d;
reg           irqarray18_eventsourceflex300_trigger_filtered;
wire          irqarray18_eventsourceflex301_status;
reg           irqarray18_eventsourceflex301_pending;
reg           irqarray18_eventsourceflex301_clear;
reg           irqarray18_eventsourceflex301_trigger_d;
reg           irqarray18_eventsourceflex301_trigger_filtered;
wire          irqarray18_eventsourceflex302_status;
reg           irqarray18_eventsourceflex302_pending;
reg           irqarray18_eventsourceflex302_clear;
reg           irqarray18_eventsourceflex302_trigger_d;
reg           irqarray18_eventsourceflex302_trigger_filtered;
wire          irqarray18_eventsourceflex303_status;
reg           irqarray18_eventsourceflex303_pending;
reg           irqarray18_eventsourceflex303_clear;
reg           irqarray18_eventsourceflex303_trigger_d;
reg           irqarray18_eventsourceflex303_trigger_filtered;
wire          irqarray18_pioirq0_dupe0;
wire          irqarray18_pioirq1_dupe0;
wire          irqarray18_pioirq2_dupe0;
wire          irqarray18_pioirq3_dupe0;
wire          irqarray18_i2c2_rx_dupe0;
wire          irqarray18_i2c2_tx_dupe0;
wire          irqarray18_i2c2_cmd_dupe0;
wire          irqarray18_i2c2_eot_dupe0;
wire          irqarray18_i2c0_nack_dupe0;
wire          irqarray18_i2c1_nack_dupe0;
wire          irqarray18_i2c2_nack_dupe0;
wire          irqarray18_i2c0_err_dupe0;
wire          irqarray18_i2c1_err_dupe0;
wire          irqarray18_i2c2_err_dupe0;
wire          irqarray18_ioxirq_dupe0;
wire          irqarray18_cam_rx_dupe0;
reg    [15:0] irqarray18_status_status;
wire          irqarray18_status_we;
reg           irqarray18_status_re;
wire          irqarray18_pioirq0_dupe1;
wire          irqarray18_pioirq1_dupe1;
wire          irqarray18_pioirq2_dupe1;
wire          irqarray18_pioirq3_dupe1;
wire          irqarray18_i2c2_rx_dupe1;
wire          irqarray18_i2c2_tx_dupe1;
wire          irqarray18_i2c2_cmd_dupe1;
wire          irqarray18_i2c2_eot_dupe1;
wire          irqarray18_i2c0_nack_dupe1;
wire          irqarray18_i2c1_nack_dupe1;
wire          irqarray18_i2c2_nack_dupe1;
wire          irqarray18_i2c0_err_dupe1;
wire          irqarray18_i2c1_err_dupe1;
wire          irqarray18_i2c2_err_dupe1;
wire          irqarray18_ioxirq_dupe1;
wire          irqarray18_cam_rx_dupe1;
reg    [15:0] irqarray18_pending_status;
wire          irqarray18_pending_we;
reg           irqarray18_pending_re;
reg    [15:0] irqarray18_pending_r;
wire          irqarray18_pioirq0_dupe2;
wire          irqarray18_pioirq1_dupe2;
wire          irqarray18_pioirq2_dupe2;
wire          irqarray18_pioirq3_dupe2;
wire          irqarray18_i2c2_rx_dupe2;
wire          irqarray18_i2c2_tx_dupe2;
wire          irqarray18_i2c2_cmd_dupe2;
wire          irqarray18_i2c2_eot_dupe2;
wire          irqarray18_i2c0_nack_dupe2;
wire          irqarray18_i2c1_nack_dupe2;
wire          irqarray18_i2c2_nack_dupe2;
wire          irqarray18_i2c0_err_dupe2;
wire          irqarray18_i2c1_err_dupe2;
wire          irqarray18_i2c2_err_dupe2;
wire          irqarray18_ioxirq_dupe2;
wire          irqarray18_cam_rx_dupe2;
reg    [15:0] irqarray18_enable_storage;
reg           irqarray18_enable_re;
wire          irqarray19_irq;
wire   [15:0] irqarray19_interrupts;
reg    [15:0] irqarray19_trigger;
reg    [15:0] irqarray19_soft_storage;
reg           irqarray19_soft_re;
wire   [15:0] irqarray19_use_edge;
reg    [15:0] irqarray19_edge_triggered_storage;
reg           irqarray19_edge_triggered_re;
wire   [15:0] irqarray19_rising;
reg    [15:0] irqarray19_polarity_storage;
reg           irqarray19_polarity_re;
wire          irqarray19_eventsourceflex304_status;
reg           irqarray19_eventsourceflex304_pending;
reg           irqarray19_eventsourceflex304_clear;
reg           irqarray19_eventsourceflex304_trigger_d;
reg           irqarray19_eventsourceflex304_trigger_filtered;
wire          irqarray19_eventsourceflex305_status;
reg           irqarray19_eventsourceflex305_pending;
reg           irqarray19_eventsourceflex305_clear;
reg           irqarray19_eventsourceflex305_trigger_d;
reg           irqarray19_eventsourceflex305_trigger_filtered;
wire          irqarray19_eventsourceflex306_status;
reg           irqarray19_eventsourceflex306_pending;
reg           irqarray19_eventsourceflex306_clear;
reg           irqarray19_eventsourceflex306_trigger_d;
reg           irqarray19_eventsourceflex306_trigger_filtered;
wire          irqarray19_eventsourceflex307_status;
reg           irqarray19_eventsourceflex307_pending;
reg           irqarray19_eventsourceflex307_clear;
reg           irqarray19_eventsourceflex307_trigger_d;
reg           irqarray19_eventsourceflex307_trigger_filtered;
wire          irqarray19_eventsourceflex308_status;
reg           irqarray19_eventsourceflex308_pending;
reg           irqarray19_eventsourceflex308_clear;
reg           irqarray19_eventsourceflex308_trigger_d;
reg           irqarray19_eventsourceflex308_trigger_filtered;
wire          irqarray19_eventsourceflex309_status;
reg           irqarray19_eventsourceflex309_pending;
reg           irqarray19_eventsourceflex309_clear;
reg           irqarray19_eventsourceflex309_trigger_d;
reg           irqarray19_eventsourceflex309_trigger_filtered;
wire          irqarray19_eventsourceflex310_status;
reg           irqarray19_eventsourceflex310_pending;
reg           irqarray19_eventsourceflex310_clear;
reg           irqarray19_eventsourceflex310_trigger_d;
reg           irqarray19_eventsourceflex310_trigger_filtered;
wire          irqarray19_eventsourceflex311_status;
reg           irqarray19_eventsourceflex311_pending;
reg           irqarray19_eventsourceflex311_clear;
reg           irqarray19_eventsourceflex311_trigger_d;
reg           irqarray19_eventsourceflex311_trigger_filtered;
wire          irqarray19_eventsourceflex312_status;
reg           irqarray19_eventsourceflex312_pending;
reg           irqarray19_eventsourceflex312_clear;
reg           irqarray19_eventsourceflex312_trigger_d;
reg           irqarray19_eventsourceflex312_trigger_filtered;
wire          irqarray19_eventsourceflex313_status;
reg           irqarray19_eventsourceflex313_pending;
reg           irqarray19_eventsourceflex313_clear;
reg           irqarray19_eventsourceflex313_trigger_d;
reg           irqarray19_eventsourceflex313_trigger_filtered;
wire          irqarray19_eventsourceflex314_status;
reg           irqarray19_eventsourceflex314_pending;
reg           irqarray19_eventsourceflex314_clear;
reg           irqarray19_eventsourceflex314_trigger_d;
reg           irqarray19_eventsourceflex314_trigger_filtered;
wire          irqarray19_eventsourceflex315_status;
reg           irqarray19_eventsourceflex315_pending;
reg           irqarray19_eventsourceflex315_clear;
reg           irqarray19_eventsourceflex315_trigger_d;
reg           irqarray19_eventsourceflex315_trigger_filtered;
wire          irqarray19_eventsourceflex316_status;
reg           irqarray19_eventsourceflex316_pending;
reg           irqarray19_eventsourceflex316_clear;
reg           irqarray19_eventsourceflex316_trigger_d;
reg           irqarray19_eventsourceflex316_trigger_filtered;
wire          irqarray19_eventsourceflex317_status;
reg           irqarray19_eventsourceflex317_pending;
reg           irqarray19_eventsourceflex317_clear;
reg           irqarray19_eventsourceflex317_trigger_d;
reg           irqarray19_eventsourceflex317_trigger_filtered;
wire          irqarray19_eventsourceflex318_status;
reg           irqarray19_eventsourceflex318_pending;
reg           irqarray19_eventsourceflex318_clear;
reg           irqarray19_eventsourceflex318_trigger_d;
reg           irqarray19_eventsourceflex318_trigger_filtered;
wire          irqarray19_eventsourceflex319_status;
reg           irqarray19_eventsourceflex319_pending;
reg           irqarray19_eventsourceflex319_clear;
reg           irqarray19_eventsourceflex319_trigger_d;
reg           irqarray19_eventsourceflex319_trigger_filtered;
wire          irqarray19_mbox_irq_available_dupe0;
wire          irqarray19_mbox_irq_abort_init_dupe0;
wire          irqarray19_mbox_irq_done_dupe0;
wire          irqarray19_mbox_irq_error_dupe0;
wire          irqarray19_pioirq0_dupe0;
wire          irqarray19_pioirq1_dupe0;
wire          irqarray19_pioirq2_dupe0;
wire          irqarray19_pioirq3_dupe0;
wire          irqarray19_sdio_rx_dupe0;
wire          irqarray19_sdio_tx_dupe0;
wire          irqarray19_sdio_eot_dupe0;
wire          irqarray19_sdio_err_dupe0;
wire          irqarray19_nc_b19s120;
wire          irqarray19_nc_b19s130;
wire          irqarray19_nc_b19s140;
wire          irqarray19_nc_b19s150;
reg    [15:0] irqarray19_status_status;
wire          irqarray19_status_we;
reg           irqarray19_status_re;
wire          irqarray19_mbox_irq_available_dupe1;
wire          irqarray19_mbox_irq_abort_init_dupe1;
wire          irqarray19_mbox_irq_done_dupe1;
wire          irqarray19_mbox_irq_error_dupe1;
wire          irqarray19_pioirq0_dupe1;
wire          irqarray19_pioirq1_dupe1;
wire          irqarray19_pioirq2_dupe1;
wire          irqarray19_pioirq3_dupe1;
wire          irqarray19_sdio_rx_dupe1;
wire          irqarray19_sdio_tx_dupe1;
wire          irqarray19_sdio_eot_dupe1;
wire          irqarray19_sdio_err_dupe1;
wire          irqarray19_nc_b19s121;
wire          irqarray19_nc_b19s131;
wire          irqarray19_nc_b19s141;
wire          irqarray19_nc_b19s151;
reg    [15:0] irqarray19_pending_status;
wire          irqarray19_pending_we;
reg           irqarray19_pending_re;
reg    [15:0] irqarray19_pending_r;
wire          irqarray19_mbox_irq_available_dupe2;
wire          irqarray19_mbox_irq_abort_init_dupe2;
wire          irqarray19_mbox_irq_done_dupe2;
wire          irqarray19_mbox_irq_error_dupe2;
wire          irqarray19_pioirq0_dupe2;
wire          irqarray19_pioirq1_dupe2;
wire          irqarray19_pioirq2_dupe2;
wire          irqarray19_pioirq3_dupe2;
wire          irqarray19_sdio_rx_dupe2;
wire          irqarray19_sdio_tx_dupe2;
wire          irqarray19_sdio_eot_dupe2;
wire          irqarray19_sdio_err_dupe2;
wire          irqarray19_nc_b19s122;
wire          irqarray19_nc_b19s132;
wire          irqarray19_nc_b19s142;
wire          irqarray19_nc_b19s152;
reg    [15:0] irqarray19_enable_storage;
reg           irqarray19_enable_re;
wire   [31:0] ticktimer_clkspertick;
reg    [31:0] ticktimer_prescaler;
reg    [63:0] ticktimer_timer0;
wire          ticktimer_pause0;
wire          ticktimer_pause1;
wire          ticktimer_load;
wire          ticktimer_load_xfer_i;
wire          ticktimer_load_xfer_o;
wire          ticktimer_load_xfer_ps_i;
wire          ticktimer_load_xfer_ps_o;
reg           ticktimer_load_xfer_ps_toggle_i;
wire          ticktimer_load_xfer_ps_toggle_o;
reg           ticktimer_load_xfer_ps_toggle_o_r;
wire          ticktimer_load_xfer_ps_ack_i;
wire          ticktimer_load_xfer_ps_ack_o;
reg           ticktimer_load_xfer_ps_ack_toggle_i;
wire          ticktimer_load_xfer_ps_ack_toggle_o;
reg           ticktimer_load_xfer_ps_ack_toggle_o_r;
reg           ticktimer_load_xfer_blind;
wire          ticktimer_paused0;
reg           ticktimer_paused1;
wire   [63:0] ticktimer_timer1;
wire   [63:0] ticktimer_timer_sync_i;
reg    [63:0] ticktimer_timer_sync_o;
reg           ticktimer_timer_sync_starter;
wire          ticktimer_timer_sync_ping_i;
wire          ticktimer_timer_sync_ping_o0;
reg           ticktimer_timer_sync_ping_toggle_i;
wire          ticktimer_timer_sync_ping_toggle_o;
reg           ticktimer_timer_sync_ping_toggle_o_r;
reg           ticktimer_timer_sync_ping_o1;
wire          ticktimer_timer_sync_pong_i;
wire          ticktimer_timer_sync_pong_o;
reg           ticktimer_timer_sync_pong_toggle_i;
wire          ticktimer_timer_sync_pong_toggle_o;
reg           ticktimer_timer_sync_pong_toggle_o_r;
wire          ticktimer_timer_sync_wait;
wire          ticktimer_timer_sync_done;
reg     [7:0] ticktimer_timer_sync_count;
reg    [63:0] ticktimer_timer_sync_ibuffer;
wire   [63:0] ticktimer_timer_sync_obuffer;
wire   [63:0] ticktimer_resume_time;
wire   [63:0] ticktimer_resume_sync_i;
reg    [63:0] ticktimer_resume_sync_o;
reg           ticktimer_resume_sync_starter;
wire          ticktimer_resume_sync_ping_i;
wire          ticktimer_resume_sync_ping_o0;
reg           ticktimer_resume_sync_ping_toggle_i;
wire          ticktimer_resume_sync_ping_toggle_o;
reg           ticktimer_resume_sync_ping_toggle_o_r;
reg           ticktimer_resume_sync_ping_o1;
wire          ticktimer_resume_sync_pong_i;
wire          ticktimer_resume_sync_pong_o;
reg           ticktimer_resume_sync_pong_toggle_i;
wire          ticktimer_resume_sync_pong_toggle_o;
reg           ticktimer_resume_sync_pong_toggle_o_r;
wire          ticktimer_resume_sync_wait;
wire          ticktimer_resume_sync_done;
reg     [7:0] ticktimer_resume_sync_count;
reg    [63:0] ticktimer_resume_sync_ibuffer;
wire   [63:0] ticktimer_resume_sync_obuffer;
reg           ticktimer_reset;
reg           ticktimer_control_storage;
reg           ticktimer_control_re;
wire   [63:0] ticktimer_time_status;
wire          ticktimer_time_we;
reg           ticktimer_time_re;
wire          ticktimer_reset_xfer_i;
wire          ticktimer_reset_xfer_o;
wire          ticktimer_reset_xfer_ps_i;
wire          ticktimer_reset_xfer_ps_o;
reg           ticktimer_reset_xfer_ps_toggle_i;
wire          ticktimer_reset_xfer_ps_toggle_o;
reg           ticktimer_reset_xfer_ps_toggle_o_r;
wire          ticktimer_reset_xfer_ps_ack_i;
wire          ticktimer_reset_xfer_ps_ack_o;
reg           ticktimer_reset_xfer_ps_ack_toggle_i;
wire          ticktimer_reset_xfer_ps_ack_toggle_o;
reg           ticktimer_reset_xfer_ps_ack_toggle_o_r;
reg           ticktimer_reset_xfer_blind;
reg    [63:0] ticktimer_msleep_target_storage;
reg           ticktimer_msleep_target_re;
wire          ticktimer_irq;
wire          ticktimer_alarm_status;
wire          ticktimer_alarm_pending;
wire          ticktimer_alarm_trigger0;
reg           ticktimer_alarm_clear;
reg           ticktimer_alarm_trigger1;
wire          ticktimer_alarm0;
wire          ticktimer_status_status;
wire          ticktimer_status_we;
reg           ticktimer_status_re;
wire          ticktimer_alarm1;
wire          ticktimer_pending_status;
wire          ticktimer_pending_we;
reg           ticktimer_pending_re;
reg           ticktimer_pending_r;
wire          ticktimer_alarm2;
reg           ticktimer_enable_storage;
reg           ticktimer_enable_re;
wire          ticktimer_ping_i;
wire          ticktimer_ping_o;
wire          ticktimer_ping_ps_i;
wire          ticktimer_ping_ps_o;
reg           ticktimer_ping_ps_toggle_i;
wire          ticktimer_ping_ps_toggle_o;
reg           ticktimer_ping_ps_toggle_o_r;
wire          ticktimer_ping_ps_ack_i;
wire          ticktimer_ping_ps_ack_o;
reg           ticktimer_ping_ps_ack_toggle_i;
wire          ticktimer_ping_ps_ack_toggle_o;
reg           ticktimer_ping_ps_ack_toggle_o_r;
reg           ticktimer_ping_blind;
wire          ticktimer_pong_i;
wire          ticktimer_pong_o;
wire          ticktimer_pong_ps_i;
wire          ticktimer_pong_ps_o;
reg           ticktimer_pong_ps_toggle_i;
wire          ticktimer_pong_ps_toggle_o;
reg           ticktimer_pong_ps_toggle_o_r;
wire          ticktimer_pong_ps_ack_i;
wire          ticktimer_pong_ps_ack_o;
reg           ticktimer_pong_ps_ack_toggle_i;
wire          ticktimer_pong_ps_ack_toggle_o;
reg           ticktimer_pong_ps_ack_toggle_o_r;
reg           ticktimer_pong_blind;
reg           ticktimer_lockout_alarm;
reg           ticktimer_alarm3;
wire   [63:0] ticktimer_target_xfer_i;
reg    [63:0] ticktimer_target_xfer_o;
reg           ticktimer_target_xfer_starter;
wire          ticktimer_target_xfer_ping_i;
wire          ticktimer_target_xfer_ping_o0;
reg           ticktimer_target_xfer_ping_toggle_i;
wire          ticktimer_target_xfer_ping_toggle_o;
reg           ticktimer_target_xfer_ping_toggle_o_r;
reg           ticktimer_target_xfer_ping_o1;
wire          ticktimer_target_xfer_pong_i;
wire          ticktimer_target_xfer_pong_o;
reg           ticktimer_target_xfer_pong_toggle_i;
wire          ticktimer_target_xfer_pong_toggle_o;
reg           ticktimer_target_xfer_pong_toggle_o_r;
wire          ticktimer_target_xfer_wait;
wire          ticktimer_target_xfer_done;
reg     [7:0] ticktimer_target_xfer_count;
reg    [63:0] ticktimer_target_xfer_ibuffer;
wire   [63:0] ticktimer_target_xfer_obuffer;
wire          ticktimer_alarm_always_on;
reg    [31:0] ticktimer_clocks_per_tick_storage;
reg           ticktimer_clocks_per_tick_re;
wire   [31:0] d11ctime_count;
reg    [31:0] d11ctime_control_storage;
reg           d11ctime_control_re;
wire          d11ctime_beat;
wire          d11ctime_heartbeat_status;
wire          d11ctime_heartbeat_we;
reg           d11ctime_heartbeat_re;
reg    [31:0] d11ctime_counter;
reg           d11ctime_heartbeat;
wire          susres_pause;
reg           susres_load;
reg     [1:0] susres_control_storage;
reg           susres_control_re;
reg    [63:0] susres_resume_time_storage;
reg           susres_resume_time_re;
wire   [63:0] susres_time_status;
wire          susres_time_we;
reg           susres_time_re;
wire          susres_paused;
wire          susres_status_status0;
wire          susres_status_we0;
reg           susres_status_re0;
wire          susres_resume0;
wire          susres_was_forced;
reg     [1:0] susres_state_storage;
reg           susres_state_re;
wire          susres_resume1;
reg           susres_interrupt;
reg           susres_interrupt_storage;
reg           susres_interrupt_re;
wire          susres_irq;
wire          susres_soft_int_status;
reg           susres_soft_int_pending;
wire          susres_soft_int_trigger;
reg           susres_soft_int_clear;
reg           susres_soft_int_trigger_d;
reg           susres_kernel_resume_interrupt;
wire          susres_soft_int0;
wire          susres_status_status1;
wire          susres_status_we1;
reg           susres_status_re1;
wire          susres_soft_int1;
wire          susres_pending_status;
wire          susres_pending_we;
reg           susres_pending_re;
reg           susres_pending_r;
wire          susres_soft_int2;
reg           susres_enable_storage;
reg           susres_enable_re;
wire          mailbox_cmatpg;
wire          mailbox_cmbist;
wire    [2:0] mailbox_vexsramtrm;
wire   [31:0] mailbox_w_dat;
wire          mailbox_w_valid;
wire          mailbox_w_ready;
wire          mailbox_w_done;
wire   [31:0] mailbox_r_dat;
wire          mailbox_r_valid;
wire          mailbox_r_ready;
wire          mailbox_r_done;
reg           mailbox_w_abort;
wire          mailbox_r_abort;
wire          mailbox_reset_n;
reg    [31:0] mailbox_wdata_storage;
reg           mailbox_wdata_re;
wire   [31:0] mailbox_rdata_status;
wire          mailbox_rdata_we;
reg           mailbox_rdata_re;
wire          mailbox_irq;
wire          mailbox_available_status;
reg           mailbox_available_pending;
wire          mailbox_available_trigger;
reg           mailbox_available_clear;
wire          mailbox_abort_init_status;
reg           mailbox_abort_init_pending;
reg           mailbox_abort_init_trigger;
reg           mailbox_abort_init_clear;
reg           mailbox_abort_init_trigger_d;
wire          mailbox_abort_done_status;
reg           mailbox_abort_done_pending;
reg           mailbox_abort_done_trigger;
reg           mailbox_abort_done_clear;
reg           mailbox_abort_done_trigger_d;
wire          mailbox_error_status;
reg           mailbox_error_pending;
wire          mailbox_error_trigger;
reg           mailbox_error_clear;
reg           mailbox_error_trigger_d;
wire          mailbox_available0;
wire          mailbox_abort_init0;
wire          mailbox_abort_done0;
wire          mailbox_error0;
reg     [3:0] mailbox_status_status0;
wire          mailbox_status_we0;
reg           mailbox_status_re0;
wire          mailbox_available1;
wire          mailbox_abort_init1;
wire          mailbox_abort_done1;
wire          mailbox_error1;
reg     [3:0] mailbox_pending_status;
wire          mailbox_pending_we;
reg           mailbox_pending_re;
reg     [3:0] mailbox_pending_r;
wire          mailbox_available2;
wire          mailbox_abort_init2;
wire          mailbox_abort_done2;
wire          mailbox_error2;
reg     [3:0] mailbox_enable_storage;
reg           mailbox_enable_re;
wire   [10:0] mailbox_rx_words;
wire   [10:0] mailbox_tx_words;
wire          mailbox_abort_in_progress0;
wire          mailbox_abort_ack0;
wire          mailbox_tx_err;
wire          mailbox_rx_err;
reg    [25:0] mailbox_status_status1;
wire          mailbox_status_we1;
reg           mailbox_status_re1;
reg           mailbox_abort;
reg           mailbox_control_storage;
reg           mailbox_control_re;
reg           mailbox_done;
reg           mailbox_done_storage;
reg           mailbox_done_re;
wire          mailbox_loopback;
reg           mailbox_loopback_storage;
reg           mailbox_loopback_re;
reg           mailbox_abort_in_progress1;
reg           mailbox_abort_ack1;
reg           mailbox_w_over_flag;
reg           mailbox_w_over_bit;
wire          mailbox_w_over_clear;
wire          mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_re;
reg           mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_readable;
wire          mailbox_syncfifobufferedmacro0_cmbist;
wire          mailbox_syncfifobufferedmacro0_cmatpg;
wire    [2:0] mailbox_syncfifobufferedmacro0_vexsramtrm;
reg           mailbox_syncfifobufferedmacro0_fifo_we;
wire          mailbox_syncfifobufferedmacro0_fifo_writable;
wire          mailbox_syncfifobufferedmacro0_fifo_re;
wire          mailbox_syncfifobufferedmacro0_fifo_readable;
wire   [31:0] mailbox_syncfifobufferedmacro0_fifo_din;
wire   [31:0] mailbox_syncfifobufferedmacro0_fifo_dout;
wire          mailbox_syncfifobufferedmacro0_fifo_cmbist;
wire          mailbox_syncfifobufferedmacro0_fifo_cmatpg;
wire    [2:0] mailbox_syncfifobufferedmacro0_fifo_vexsramtrm;
reg    [10:0] mailbox_syncfifobufferedmacro0_fifo_level;
reg     [9:0] mailbox_syncfifobufferedmacro0_fifo_produce;
reg     [9:0] mailbox_syncfifobufferedmacro0_fifo_consume;
reg     [9:0] mailbox_syncfifobufferedmacro0_fifo_wrport_adr;
wire   [31:0] mailbox_syncfifobufferedmacro0_fifo_wrport_dat_w;
wire          mailbox_syncfifobufferedmacro0_fifo_wrport_we;
wire    [9:0] mailbox_syncfifobufferedmacro0_fifo_rdport_adr;
wire          mailbox_syncfifobufferedmacro0_fifo_rdport_re;
wire   [31:0] mailbox_syncfifobufferedmacro0_fifo_rdport_dat_r;
wire          mailbox_syncfifobufferedmacro0_fifo_do_read;
wire   [10:0] mailbox_syncfifobufferedmacro0_level;
wire          mailbox_w_fifo_reset_sys;
reg           mailbox_r_over_flag;
reg           mailbox_r_over_bit;
wire          mailbox_r_over_clear;
reg           mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_re;
reg           mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_readable;
wire          mailbox_syncfifobufferedmacro1_cmbist;
wire          mailbox_syncfifobufferedmacro1_cmatpg;
wire    [2:0] mailbox_syncfifobufferedmacro1_vexsramtrm;
wire          mailbox_syncfifobufferedmacro1_fifo_we;
wire          mailbox_syncfifobufferedmacro1_fifo_writable;
wire          mailbox_syncfifobufferedmacro1_fifo_re;
wire          mailbox_syncfifobufferedmacro1_fifo_readable;
wire   [31:0] mailbox_syncfifobufferedmacro1_fifo_din;
wire   [31:0] mailbox_syncfifobufferedmacro1_fifo_dout;
wire          mailbox_syncfifobufferedmacro1_fifo_cmbist;
wire          mailbox_syncfifobufferedmacro1_fifo_cmatpg;
wire    [2:0] mailbox_syncfifobufferedmacro1_fifo_vexsramtrm;
reg    [10:0] mailbox_syncfifobufferedmacro1_fifo_level;
reg     [9:0] mailbox_syncfifobufferedmacro1_fifo_produce;
reg     [9:0] mailbox_syncfifobufferedmacro1_fifo_consume;
reg     [9:0] mailbox_syncfifobufferedmacro1_fifo_wrport_adr;
wire   [31:0] mailbox_syncfifobufferedmacro1_fifo_wrport_dat_w;
wire          mailbox_syncfifobufferedmacro1_fifo_wrport_we;
wire    [9:0] mailbox_syncfifobufferedmacro1_fifo_rdport_adr;
wire          mailbox_syncfifobufferedmacro1_fifo_rdport_re;
wire   [31:0] mailbox_syncfifobufferedmacro1_fifo_rdport_dat_r;
wire          mailbox_syncfifobufferedmacro1_fifo_do_read;
wire   [10:0] mailbox_syncfifobufferedmacro1_level;
wire          mailbox_r_fifo_reset_sys;
wire   [31:0] mb_client_w_dat;
wire          mb_client_w_valid;
wire          mb_client_w_ready;
wire          mb_client_w_done;
wire   [31:0] mb_client_r_dat;
wire          mb_client_r_valid;
wire          mb_client_r_ready;
wire          mb_client_r_done;
reg           mb_client_w_abort;
wire          mb_client_r_abort;
reg           mb_client_reset_n;
reg    [31:0] mb_client_wdata_storage;
reg           mb_client_wdata_re;
wire   [31:0] mb_client_rdata_status;
wire          mb_client_rdata_we;
reg           mb_client_rdata_re;
wire          mb_client_rx_avail;
wire          mb_client_tx_free;
wire          mb_client_abort_in_progress0;
wire          mb_client_abort_ack0;
reg           mb_client_tx_err;
reg           mb_client_rx_err;
reg     [5:0] mb_client_status_status0;
wire          mb_client_status_we0;
reg           mb_client_status_re0;
wire          mb_client_irq;
wire          mb_client_available_status;
reg           mb_client_available_pending;
wire          mb_client_available_trigger;
reg           mb_client_available_clear;
wire          mb_client_abort_init_status;
reg           mb_client_abort_init_pending;
reg           mb_client_abort_init_trigger;
reg           mb_client_abort_init_clear;
reg           mb_client_abort_init_trigger_d;
wire          mb_client_abort_done_status;
reg           mb_client_abort_done_pending;
reg           mb_client_abort_done_trigger;
reg           mb_client_abort_done_clear;
reg           mb_client_abort_done_trigger_d;
wire          mb_client_error_status;
reg           mb_client_error_pending;
wire          mb_client_error_trigger;
reg           mb_client_error_clear;
reg           mb_client_error_trigger_d;
wire          mb_client_available0;
wire          mb_client_abort_init0;
wire          mb_client_abort_done0;
wire          mb_client_error0;
reg     [3:0] mb_client_status_status1;
wire          mb_client_status_we1;
reg           mb_client_status_re1;
wire          mb_client_available1;
wire          mb_client_abort_init1;
wire          mb_client_abort_done1;
wire          mb_client_error1;
reg     [3:0] mb_client_pending_status;
wire          mb_client_pending_we;
reg           mb_client_pending_re;
reg     [3:0] mb_client_pending_r;
wire          mb_client_available2;
wire          mb_client_abort_init2;
wire          mb_client_abort_done2;
wire          mb_client_error2;
reg     [3:0] mb_client_enable_storage;
reg           mb_client_enable_re;
reg           mb_client_abort;
reg           mb_client_control_storage;
reg           mb_client_control_re;
reg           mb_client_done;
reg           mb_client_done_storage;
reg           mb_client_done_re;
reg           mb_client_abort_in_progress1;
reg           mb_client_abort_ack1;
reg           mb_client_w_pending;
wire          loopback;
wire   [31:0] w_dat;
wire          w_valid;
reg           w_ready;
wire          w_done;
reg    [31:0] r_dat;
reg           r_valid;
wire          r_ready;
reg           r_done;
wire          w_abort;
reg           r_abort;
reg    [31:0] csr_wtest_storage;
reg           csr_wtest_re;
wire   [31:0] csr_rtest_status;
wire          csr_rtest_we;
reg           csr_rtest_re;
reg    [15:0] cramsoc_adr;
wire          cramsoc_we;
wire   [31:0] cramsoc_dat_w;
wire   [31:0] cramsoc_dat_r;
wire          cramsoc_re;
wire          cramsoc_aw_valid;
wire          cramsoc_aw_ready;
wire          cramsoc_aw_first;
wire          cramsoc_aw_last;
wire   [31:0] cramsoc_aw_payload_addr;
wire    [2:0] cramsoc_aw_payload_prot;
wire          cramsoc_w_valid;
wire          cramsoc_w_ready;
wire          cramsoc_w_first;
wire          cramsoc_w_last;
wire   [31:0] cramsoc_w_payload_data;
wire    [3:0] cramsoc_w_payload_strb;
wire          cramsoc_b_valid;
wire          cramsoc_b_ready;
reg           cramsoc_b_first;
reg           cramsoc_b_last;
reg     [1:0] cramsoc_b_payload_resp;
wire          cramsoc_ar_valid;
wire          cramsoc_ar_ready;
wire          cramsoc_ar_first;
wire          cramsoc_ar_last;
wire   [31:0] cramsoc_ar_payload_addr;
wire    [2:0] cramsoc_ar_payload_prot;
wire          cramsoc_r_valid;
wire          cramsoc_r_ready;
reg           cramsoc_r_first;
reg           cramsoc_r_last;
reg     [1:0] cramsoc_r_payload_resp;
reg    [31:0] cramsoc_r_payload_data;
reg           cramsoc_do_read;
reg           cramsoc_do_write;
reg           cramsoc_last_was_read;
reg           cramsoc_nocomb_axl_r_valid;
reg           cramsoc_nocomb_axl_w_ready;
reg           cramsoc_nocomb_axl_aw_ready;
reg           cramsoc_nocomb_axl_ar_ready;
reg           cramsoc_nocomb_axl_b_valid;
wire          socbushandler_aw_valid;
reg           socbushandler_aw_ready;
wire          socbushandler_aw_first;
wire          socbushandler_aw_last;
wire   [31:0] socbushandler_aw_payload_addr;
wire    [2:0] socbushandler_aw_payload_prot;
wire          socbushandler_w_valid;
reg           socbushandler_w_ready;
wire          socbushandler_w_first;
wire          socbushandler_w_last;
wire   [31:0] socbushandler_w_payload_data;
wire    [3:0] socbushandler_w_payload_strb;
reg           socbushandler_b_valid;
wire          socbushandler_b_ready;
wire          socbushandler_b_first;
wire          socbushandler_b_last;
wire    [1:0] socbushandler_b_payload_resp;
wire          socbushandler_ar_valid;
reg           socbushandler_ar_ready;
wire          socbushandler_ar_first;
wire          socbushandler_ar_last;
wire   [31:0] socbushandler_ar_payload_addr;
wire    [2:0] socbushandler_ar_payload_prot;
reg           socbushandler_r_valid;
wire          socbushandler_r_ready;
wire          socbushandler_r_first;
wire          socbushandler_r_last;
wire    [1:0] socbushandler_r_payload_resp;
wire   [31:0] socbushandler_r_payload_data;
wire          socbushandler_slave_sel_dec0;
wire          socbushandler_slave_sel_dec1;
reg           socbushandler_slave_sel_reg0;
reg           socbushandler_slave_sel_reg1;
reg           socbushandler_slave_sel0;
reg           socbushandler_slave_sel1;
reg     [7:0] socbushandler_axiliterequestcounter0_counter;
wire          socbushandler_axiliterequestcounter0_full;
wire          socbushandler_axiliterequestcounter0_empty;
wire          socbushandler_axiliterequestcounter0_stall;
reg     [7:0] socbushandler_axiliterequestcounter1_counter;
wire          socbushandler_axiliterequestcounter1_full;
wire          socbushandler_axiliterequestcounter1_empty;
wire          socbushandler_axiliterequestcounter1_stall;
wire          socbushandler_rr_write_request;
wire          socbushandler_rr_write_grant;
wire          socbushandler_rr_write_ce;
wire          socbushandler_rr_read_request;
wire          socbushandler_rr_read_grant;
wire          socbushandler_rr_read_ce;
reg     [7:0] socbushandler_wr_lock_counter;
wire          socbushandler_wr_lock_full;
wire          socbushandler_wr_lock_empty;
wire          socbushandler_wr_lock_stall;
reg     [7:0] socbushandler_rd_lock_counter;
wire          socbushandler_rd_lock_full;
wire          socbushandler_rd_lock_empty;
wire          socbushandler_rd_lock_stall;
wire   [15:0] interface0_bank_bus_adr;
wire          interface0_bank_bus_we;
wire   [31:0] interface0_bank_bus_dat_w;
reg    [31:0] interface0_bank_bus_dat_r;
wire          interface0_bank_bus_re;
reg           csrbank0_control0_re;
wire    [1:0] csrbank0_control0_r;
reg           csrbank0_control0_we;
wire    [1:0] csrbank0_control0_w;
reg           csrbank0_status_re;
wire    [8:0] csrbank0_status_r;
reg           csrbank0_status_we;
wire    [8:0] csrbank0_status_w;
reg           csrbank0_map_lo0_re;
wire   [31:0] csrbank0_map_lo0_r;
reg           csrbank0_map_lo0_we;
wire   [31:0] csrbank0_map_lo0_w;
reg           csrbank0_map_hi0_re;
wire   [31:0] csrbank0_map_hi0_r;
reg           csrbank0_map_hi0_we;
wire   [31:0] csrbank0_map_hi0_w;
reg           csrbank0_uservalue0_re;
wire   [17:0] csrbank0_uservalue0_r;
reg           csrbank0_uservalue0_we;
wire   [17:0] csrbank0_uservalue0_w;
reg           csrbank0_protect0_re;
wire          csrbank0_protect0_r;
reg           csrbank0_protect0_we;
wire          csrbank0_protect0_w;
wire          csrbank0_sel;
wire          csrbank0_re;
wire   [15:0] interface1_bank_bus_adr;
wire          interface1_bank_bus_we;
wire   [31:0] interface1_bank_bus_dat_w;
reg    [31:0] interface1_bank_bus_dat_r;
wire          interface1_bank_bus_re;
reg           csrbank1_wtest0_re;
wire   [31:0] csrbank1_wtest0_r;
reg           csrbank1_wtest0_we;
wire   [31:0] csrbank1_wtest0_w;
reg           csrbank1_rtest_re;
wire   [31:0] csrbank1_rtest_r;
reg           csrbank1_rtest_we;
wire   [31:0] csrbank1_rtest_w;
wire          csrbank1_sel;
wire          csrbank1_re;
wire   [15:0] interface2_bank_bus_adr;
wire          interface2_bank_bus_we;
wire   [31:0] interface2_bank_bus_dat_w;
reg    [31:0] interface2_bank_bus_dat_r;
wire          interface2_bank_bus_re;
reg           csrbank2_control0_re;
wire   [31:0] csrbank2_control0_r;
reg           csrbank2_control0_we;
wire   [31:0] csrbank2_control0_w;
reg           csrbank2_heartbeat_re;
wire          csrbank2_heartbeat_r;
reg           csrbank2_heartbeat_we;
wire          csrbank2_heartbeat_w;
wire          csrbank2_sel;
wire          csrbank2_re;
wire   [15:0] interface3_bank_bus_adr;
wire          interface3_bank_bus_we;
wire   [31:0] interface3_bank_bus_dat_w;
reg    [31:0] interface3_bank_bus_dat_r;
wire          interface3_bank_bus_re;
reg           csrbank3_ev_soft0_re;
wire   [15:0] csrbank3_ev_soft0_r;
reg           csrbank3_ev_soft0_we;
wire   [15:0] csrbank3_ev_soft0_w;
reg           csrbank3_ev_edge_triggered0_re;
wire   [15:0] csrbank3_ev_edge_triggered0_r;
reg           csrbank3_ev_edge_triggered0_we;
wire   [15:0] csrbank3_ev_edge_triggered0_w;
reg           csrbank3_ev_polarity0_re;
wire   [15:0] csrbank3_ev_polarity0_r;
reg           csrbank3_ev_polarity0_we;
wire   [15:0] csrbank3_ev_polarity0_w;
reg           csrbank3_ev_status_re;
wire   [15:0] csrbank3_ev_status_r;
reg           csrbank3_ev_status_we;
wire   [15:0] csrbank3_ev_status_w;
reg           csrbank3_ev_pending_re;
wire   [15:0] csrbank3_ev_pending_r;
reg           csrbank3_ev_pending_we;
wire   [15:0] csrbank3_ev_pending_w;
reg           csrbank3_ev_enable0_re;
wire   [15:0] csrbank3_ev_enable0_r;
reg           csrbank3_ev_enable0_we;
wire   [15:0] csrbank3_ev_enable0_w;
wire          csrbank3_sel;
wire          csrbank3_re;
wire   [15:0] interface4_bank_bus_adr;
wire          interface4_bank_bus_we;
wire   [31:0] interface4_bank_bus_dat_w;
reg    [31:0] interface4_bank_bus_dat_r;
wire          interface4_bank_bus_re;
reg           csrbank4_ev_soft0_re;
wire   [15:0] csrbank4_ev_soft0_r;
reg           csrbank4_ev_soft0_we;
wire   [15:0] csrbank4_ev_soft0_w;
reg           csrbank4_ev_edge_triggered0_re;
wire   [15:0] csrbank4_ev_edge_triggered0_r;
reg           csrbank4_ev_edge_triggered0_we;
wire   [15:0] csrbank4_ev_edge_triggered0_w;
reg           csrbank4_ev_polarity0_re;
wire   [15:0] csrbank4_ev_polarity0_r;
reg           csrbank4_ev_polarity0_we;
wire   [15:0] csrbank4_ev_polarity0_w;
reg           csrbank4_ev_status_re;
wire   [15:0] csrbank4_ev_status_r;
reg           csrbank4_ev_status_we;
wire   [15:0] csrbank4_ev_status_w;
reg           csrbank4_ev_pending_re;
wire   [15:0] csrbank4_ev_pending_r;
reg           csrbank4_ev_pending_we;
wire   [15:0] csrbank4_ev_pending_w;
reg           csrbank4_ev_enable0_re;
wire   [15:0] csrbank4_ev_enable0_r;
reg           csrbank4_ev_enable0_we;
wire   [15:0] csrbank4_ev_enable0_w;
wire          csrbank4_sel;
wire          csrbank4_re;
wire   [15:0] interface5_bank_bus_adr;
wire          interface5_bank_bus_we;
wire   [31:0] interface5_bank_bus_dat_w;
reg    [31:0] interface5_bank_bus_dat_r;
wire          interface5_bank_bus_re;
reg           csrbank5_ev_soft0_re;
wire   [15:0] csrbank5_ev_soft0_r;
reg           csrbank5_ev_soft0_we;
wire   [15:0] csrbank5_ev_soft0_w;
reg           csrbank5_ev_edge_triggered0_re;
wire   [15:0] csrbank5_ev_edge_triggered0_r;
reg           csrbank5_ev_edge_triggered0_we;
wire   [15:0] csrbank5_ev_edge_triggered0_w;
reg           csrbank5_ev_polarity0_re;
wire   [15:0] csrbank5_ev_polarity0_r;
reg           csrbank5_ev_polarity0_we;
wire   [15:0] csrbank5_ev_polarity0_w;
reg           csrbank5_ev_status_re;
wire   [15:0] csrbank5_ev_status_r;
reg           csrbank5_ev_status_we;
wire   [15:0] csrbank5_ev_status_w;
reg           csrbank5_ev_pending_re;
wire   [15:0] csrbank5_ev_pending_r;
reg           csrbank5_ev_pending_we;
wire   [15:0] csrbank5_ev_pending_w;
reg           csrbank5_ev_enable0_re;
wire   [15:0] csrbank5_ev_enable0_r;
reg           csrbank5_ev_enable0_we;
wire   [15:0] csrbank5_ev_enable0_w;
wire          csrbank5_sel;
wire          csrbank5_re;
wire   [15:0] interface6_bank_bus_adr;
wire          interface6_bank_bus_we;
wire   [31:0] interface6_bank_bus_dat_w;
reg    [31:0] interface6_bank_bus_dat_r;
wire          interface6_bank_bus_re;
reg           csrbank6_ev_soft0_re;
wire   [15:0] csrbank6_ev_soft0_r;
reg           csrbank6_ev_soft0_we;
wire   [15:0] csrbank6_ev_soft0_w;
reg           csrbank6_ev_edge_triggered0_re;
wire   [15:0] csrbank6_ev_edge_triggered0_r;
reg           csrbank6_ev_edge_triggered0_we;
wire   [15:0] csrbank6_ev_edge_triggered0_w;
reg           csrbank6_ev_polarity0_re;
wire   [15:0] csrbank6_ev_polarity0_r;
reg           csrbank6_ev_polarity0_we;
wire   [15:0] csrbank6_ev_polarity0_w;
reg           csrbank6_ev_status_re;
wire   [15:0] csrbank6_ev_status_r;
reg           csrbank6_ev_status_we;
wire   [15:0] csrbank6_ev_status_w;
reg           csrbank6_ev_pending_re;
wire   [15:0] csrbank6_ev_pending_r;
reg           csrbank6_ev_pending_we;
wire   [15:0] csrbank6_ev_pending_w;
reg           csrbank6_ev_enable0_re;
wire   [15:0] csrbank6_ev_enable0_r;
reg           csrbank6_ev_enable0_we;
wire   [15:0] csrbank6_ev_enable0_w;
wire          csrbank6_sel;
wire          csrbank6_re;
wire   [15:0] interface7_bank_bus_adr;
wire          interface7_bank_bus_we;
wire   [31:0] interface7_bank_bus_dat_w;
reg    [31:0] interface7_bank_bus_dat_r;
wire          interface7_bank_bus_re;
reg           csrbank7_ev_soft0_re;
wire   [15:0] csrbank7_ev_soft0_r;
reg           csrbank7_ev_soft0_we;
wire   [15:0] csrbank7_ev_soft0_w;
reg           csrbank7_ev_edge_triggered0_re;
wire   [15:0] csrbank7_ev_edge_triggered0_r;
reg           csrbank7_ev_edge_triggered0_we;
wire   [15:0] csrbank7_ev_edge_triggered0_w;
reg           csrbank7_ev_polarity0_re;
wire   [15:0] csrbank7_ev_polarity0_r;
reg           csrbank7_ev_polarity0_we;
wire   [15:0] csrbank7_ev_polarity0_w;
reg           csrbank7_ev_status_re;
wire   [15:0] csrbank7_ev_status_r;
reg           csrbank7_ev_status_we;
wire   [15:0] csrbank7_ev_status_w;
reg           csrbank7_ev_pending_re;
wire   [15:0] csrbank7_ev_pending_r;
reg           csrbank7_ev_pending_we;
wire   [15:0] csrbank7_ev_pending_w;
reg           csrbank7_ev_enable0_re;
wire   [15:0] csrbank7_ev_enable0_r;
reg           csrbank7_ev_enable0_we;
wire   [15:0] csrbank7_ev_enable0_w;
wire          csrbank7_sel;
wire          csrbank7_re;
wire   [15:0] interface8_bank_bus_adr;
wire          interface8_bank_bus_we;
wire   [31:0] interface8_bank_bus_dat_w;
reg    [31:0] interface8_bank_bus_dat_r;
wire          interface8_bank_bus_re;
reg           csrbank8_ev_soft0_re;
wire   [15:0] csrbank8_ev_soft0_r;
reg           csrbank8_ev_soft0_we;
wire   [15:0] csrbank8_ev_soft0_w;
reg           csrbank8_ev_edge_triggered0_re;
wire   [15:0] csrbank8_ev_edge_triggered0_r;
reg           csrbank8_ev_edge_triggered0_we;
wire   [15:0] csrbank8_ev_edge_triggered0_w;
reg           csrbank8_ev_polarity0_re;
wire   [15:0] csrbank8_ev_polarity0_r;
reg           csrbank8_ev_polarity0_we;
wire   [15:0] csrbank8_ev_polarity0_w;
reg           csrbank8_ev_status_re;
wire   [15:0] csrbank8_ev_status_r;
reg           csrbank8_ev_status_we;
wire   [15:0] csrbank8_ev_status_w;
reg           csrbank8_ev_pending_re;
wire   [15:0] csrbank8_ev_pending_r;
reg           csrbank8_ev_pending_we;
wire   [15:0] csrbank8_ev_pending_w;
reg           csrbank8_ev_enable0_re;
wire   [15:0] csrbank8_ev_enable0_r;
reg           csrbank8_ev_enable0_we;
wire   [15:0] csrbank8_ev_enable0_w;
wire          csrbank8_sel;
wire          csrbank8_re;
wire   [15:0] interface9_bank_bus_adr;
wire          interface9_bank_bus_we;
wire   [31:0] interface9_bank_bus_dat_w;
reg    [31:0] interface9_bank_bus_dat_r;
wire          interface9_bank_bus_re;
reg           csrbank9_ev_soft0_re;
wire   [15:0] csrbank9_ev_soft0_r;
reg           csrbank9_ev_soft0_we;
wire   [15:0] csrbank9_ev_soft0_w;
reg           csrbank9_ev_edge_triggered0_re;
wire   [15:0] csrbank9_ev_edge_triggered0_r;
reg           csrbank9_ev_edge_triggered0_we;
wire   [15:0] csrbank9_ev_edge_triggered0_w;
reg           csrbank9_ev_polarity0_re;
wire   [15:0] csrbank9_ev_polarity0_r;
reg           csrbank9_ev_polarity0_we;
wire   [15:0] csrbank9_ev_polarity0_w;
reg           csrbank9_ev_status_re;
wire   [15:0] csrbank9_ev_status_r;
reg           csrbank9_ev_status_we;
wire   [15:0] csrbank9_ev_status_w;
reg           csrbank9_ev_pending_re;
wire   [15:0] csrbank9_ev_pending_r;
reg           csrbank9_ev_pending_we;
wire   [15:0] csrbank9_ev_pending_w;
reg           csrbank9_ev_enable0_re;
wire   [15:0] csrbank9_ev_enable0_r;
reg           csrbank9_ev_enable0_we;
wire   [15:0] csrbank9_ev_enable0_w;
wire          csrbank9_sel;
wire          csrbank9_re;
wire   [15:0] interface10_bank_bus_adr;
wire          interface10_bank_bus_we;
wire   [31:0] interface10_bank_bus_dat_w;
reg    [31:0] interface10_bank_bus_dat_r;
wire          interface10_bank_bus_re;
reg           csrbank10_ev_soft0_re;
wire   [15:0] csrbank10_ev_soft0_r;
reg           csrbank10_ev_soft0_we;
wire   [15:0] csrbank10_ev_soft0_w;
reg           csrbank10_ev_edge_triggered0_re;
wire   [15:0] csrbank10_ev_edge_triggered0_r;
reg           csrbank10_ev_edge_triggered0_we;
wire   [15:0] csrbank10_ev_edge_triggered0_w;
reg           csrbank10_ev_polarity0_re;
wire   [15:0] csrbank10_ev_polarity0_r;
reg           csrbank10_ev_polarity0_we;
wire   [15:0] csrbank10_ev_polarity0_w;
reg           csrbank10_ev_status_re;
wire   [15:0] csrbank10_ev_status_r;
reg           csrbank10_ev_status_we;
wire   [15:0] csrbank10_ev_status_w;
reg           csrbank10_ev_pending_re;
wire   [15:0] csrbank10_ev_pending_r;
reg           csrbank10_ev_pending_we;
wire   [15:0] csrbank10_ev_pending_w;
reg           csrbank10_ev_enable0_re;
wire   [15:0] csrbank10_ev_enable0_r;
reg           csrbank10_ev_enable0_we;
wire   [15:0] csrbank10_ev_enable0_w;
wire          csrbank10_sel;
wire          csrbank10_re;
wire   [15:0] interface11_bank_bus_adr;
wire          interface11_bank_bus_we;
wire   [31:0] interface11_bank_bus_dat_w;
reg    [31:0] interface11_bank_bus_dat_r;
wire          interface11_bank_bus_re;
reg           csrbank11_ev_soft0_re;
wire   [15:0] csrbank11_ev_soft0_r;
reg           csrbank11_ev_soft0_we;
wire   [15:0] csrbank11_ev_soft0_w;
reg           csrbank11_ev_edge_triggered0_re;
wire   [15:0] csrbank11_ev_edge_triggered0_r;
reg           csrbank11_ev_edge_triggered0_we;
wire   [15:0] csrbank11_ev_edge_triggered0_w;
reg           csrbank11_ev_polarity0_re;
wire   [15:0] csrbank11_ev_polarity0_r;
reg           csrbank11_ev_polarity0_we;
wire   [15:0] csrbank11_ev_polarity0_w;
reg           csrbank11_ev_status_re;
wire   [15:0] csrbank11_ev_status_r;
reg           csrbank11_ev_status_we;
wire   [15:0] csrbank11_ev_status_w;
reg           csrbank11_ev_pending_re;
wire   [15:0] csrbank11_ev_pending_r;
reg           csrbank11_ev_pending_we;
wire   [15:0] csrbank11_ev_pending_w;
reg           csrbank11_ev_enable0_re;
wire   [15:0] csrbank11_ev_enable0_r;
reg           csrbank11_ev_enable0_we;
wire   [15:0] csrbank11_ev_enable0_w;
wire          csrbank11_sel;
wire          csrbank11_re;
wire   [15:0] interface12_bank_bus_adr;
wire          interface12_bank_bus_we;
wire   [31:0] interface12_bank_bus_dat_w;
reg    [31:0] interface12_bank_bus_dat_r;
wire          interface12_bank_bus_re;
reg           csrbank12_ev_soft0_re;
wire   [15:0] csrbank12_ev_soft0_r;
reg           csrbank12_ev_soft0_we;
wire   [15:0] csrbank12_ev_soft0_w;
reg           csrbank12_ev_edge_triggered0_re;
wire   [15:0] csrbank12_ev_edge_triggered0_r;
reg           csrbank12_ev_edge_triggered0_we;
wire   [15:0] csrbank12_ev_edge_triggered0_w;
reg           csrbank12_ev_polarity0_re;
wire   [15:0] csrbank12_ev_polarity0_r;
reg           csrbank12_ev_polarity0_we;
wire   [15:0] csrbank12_ev_polarity0_w;
reg           csrbank12_ev_status_re;
wire   [15:0] csrbank12_ev_status_r;
reg           csrbank12_ev_status_we;
wire   [15:0] csrbank12_ev_status_w;
reg           csrbank12_ev_pending_re;
wire   [15:0] csrbank12_ev_pending_r;
reg           csrbank12_ev_pending_we;
wire   [15:0] csrbank12_ev_pending_w;
reg           csrbank12_ev_enable0_re;
wire   [15:0] csrbank12_ev_enable0_r;
reg           csrbank12_ev_enable0_we;
wire   [15:0] csrbank12_ev_enable0_w;
wire          csrbank12_sel;
wire          csrbank12_re;
wire   [15:0] interface13_bank_bus_adr;
wire          interface13_bank_bus_we;
wire   [31:0] interface13_bank_bus_dat_w;
reg    [31:0] interface13_bank_bus_dat_r;
wire          interface13_bank_bus_re;
reg           csrbank13_ev_soft0_re;
wire   [15:0] csrbank13_ev_soft0_r;
reg           csrbank13_ev_soft0_we;
wire   [15:0] csrbank13_ev_soft0_w;
reg           csrbank13_ev_edge_triggered0_re;
wire   [15:0] csrbank13_ev_edge_triggered0_r;
reg           csrbank13_ev_edge_triggered0_we;
wire   [15:0] csrbank13_ev_edge_triggered0_w;
reg           csrbank13_ev_polarity0_re;
wire   [15:0] csrbank13_ev_polarity0_r;
reg           csrbank13_ev_polarity0_we;
wire   [15:0] csrbank13_ev_polarity0_w;
reg           csrbank13_ev_status_re;
wire   [15:0] csrbank13_ev_status_r;
reg           csrbank13_ev_status_we;
wire   [15:0] csrbank13_ev_status_w;
reg           csrbank13_ev_pending_re;
wire   [15:0] csrbank13_ev_pending_r;
reg           csrbank13_ev_pending_we;
wire   [15:0] csrbank13_ev_pending_w;
reg           csrbank13_ev_enable0_re;
wire   [15:0] csrbank13_ev_enable0_r;
reg           csrbank13_ev_enable0_we;
wire   [15:0] csrbank13_ev_enable0_w;
wire          csrbank13_sel;
wire          csrbank13_re;
wire   [15:0] interface14_bank_bus_adr;
wire          interface14_bank_bus_we;
wire   [31:0] interface14_bank_bus_dat_w;
reg    [31:0] interface14_bank_bus_dat_r;
wire          interface14_bank_bus_re;
reg           csrbank14_ev_soft0_re;
wire   [15:0] csrbank14_ev_soft0_r;
reg           csrbank14_ev_soft0_we;
wire   [15:0] csrbank14_ev_soft0_w;
reg           csrbank14_ev_edge_triggered0_re;
wire   [15:0] csrbank14_ev_edge_triggered0_r;
reg           csrbank14_ev_edge_triggered0_we;
wire   [15:0] csrbank14_ev_edge_triggered0_w;
reg           csrbank14_ev_polarity0_re;
wire   [15:0] csrbank14_ev_polarity0_r;
reg           csrbank14_ev_polarity0_we;
wire   [15:0] csrbank14_ev_polarity0_w;
reg           csrbank14_ev_status_re;
wire   [15:0] csrbank14_ev_status_r;
reg           csrbank14_ev_status_we;
wire   [15:0] csrbank14_ev_status_w;
reg           csrbank14_ev_pending_re;
wire   [15:0] csrbank14_ev_pending_r;
reg           csrbank14_ev_pending_we;
wire   [15:0] csrbank14_ev_pending_w;
reg           csrbank14_ev_enable0_re;
wire   [15:0] csrbank14_ev_enable0_r;
reg           csrbank14_ev_enable0_we;
wire   [15:0] csrbank14_ev_enable0_w;
wire          csrbank14_sel;
wire          csrbank14_re;
wire   [15:0] interface15_bank_bus_adr;
wire          interface15_bank_bus_we;
wire   [31:0] interface15_bank_bus_dat_w;
reg    [31:0] interface15_bank_bus_dat_r;
wire          interface15_bank_bus_re;
reg           csrbank15_ev_soft0_re;
wire   [15:0] csrbank15_ev_soft0_r;
reg           csrbank15_ev_soft0_we;
wire   [15:0] csrbank15_ev_soft0_w;
reg           csrbank15_ev_edge_triggered0_re;
wire   [15:0] csrbank15_ev_edge_triggered0_r;
reg           csrbank15_ev_edge_triggered0_we;
wire   [15:0] csrbank15_ev_edge_triggered0_w;
reg           csrbank15_ev_polarity0_re;
wire   [15:0] csrbank15_ev_polarity0_r;
reg           csrbank15_ev_polarity0_we;
wire   [15:0] csrbank15_ev_polarity0_w;
reg           csrbank15_ev_status_re;
wire   [15:0] csrbank15_ev_status_r;
reg           csrbank15_ev_status_we;
wire   [15:0] csrbank15_ev_status_w;
reg           csrbank15_ev_pending_re;
wire   [15:0] csrbank15_ev_pending_r;
reg           csrbank15_ev_pending_we;
wire   [15:0] csrbank15_ev_pending_w;
reg           csrbank15_ev_enable0_re;
wire   [15:0] csrbank15_ev_enable0_r;
reg           csrbank15_ev_enable0_we;
wire   [15:0] csrbank15_ev_enable0_w;
wire          csrbank15_sel;
wire          csrbank15_re;
wire   [15:0] interface16_bank_bus_adr;
wire          interface16_bank_bus_we;
wire   [31:0] interface16_bank_bus_dat_w;
reg    [31:0] interface16_bank_bus_dat_r;
wire          interface16_bank_bus_re;
reg           csrbank16_ev_soft0_re;
wire   [15:0] csrbank16_ev_soft0_r;
reg           csrbank16_ev_soft0_we;
wire   [15:0] csrbank16_ev_soft0_w;
reg           csrbank16_ev_edge_triggered0_re;
wire   [15:0] csrbank16_ev_edge_triggered0_r;
reg           csrbank16_ev_edge_triggered0_we;
wire   [15:0] csrbank16_ev_edge_triggered0_w;
reg           csrbank16_ev_polarity0_re;
wire   [15:0] csrbank16_ev_polarity0_r;
reg           csrbank16_ev_polarity0_we;
wire   [15:0] csrbank16_ev_polarity0_w;
reg           csrbank16_ev_status_re;
wire   [15:0] csrbank16_ev_status_r;
reg           csrbank16_ev_status_we;
wire   [15:0] csrbank16_ev_status_w;
reg           csrbank16_ev_pending_re;
wire   [15:0] csrbank16_ev_pending_r;
reg           csrbank16_ev_pending_we;
wire   [15:0] csrbank16_ev_pending_w;
reg           csrbank16_ev_enable0_re;
wire   [15:0] csrbank16_ev_enable0_r;
reg           csrbank16_ev_enable0_we;
wire   [15:0] csrbank16_ev_enable0_w;
wire          csrbank16_sel;
wire          csrbank16_re;
wire   [15:0] interface17_bank_bus_adr;
wire          interface17_bank_bus_we;
wire   [31:0] interface17_bank_bus_dat_w;
reg    [31:0] interface17_bank_bus_dat_r;
wire          interface17_bank_bus_re;
reg           csrbank17_ev_soft0_re;
wire   [15:0] csrbank17_ev_soft0_r;
reg           csrbank17_ev_soft0_we;
wire   [15:0] csrbank17_ev_soft0_w;
reg           csrbank17_ev_edge_triggered0_re;
wire   [15:0] csrbank17_ev_edge_triggered0_r;
reg           csrbank17_ev_edge_triggered0_we;
wire   [15:0] csrbank17_ev_edge_triggered0_w;
reg           csrbank17_ev_polarity0_re;
wire   [15:0] csrbank17_ev_polarity0_r;
reg           csrbank17_ev_polarity0_we;
wire   [15:0] csrbank17_ev_polarity0_w;
reg           csrbank17_ev_status_re;
wire   [15:0] csrbank17_ev_status_r;
reg           csrbank17_ev_status_we;
wire   [15:0] csrbank17_ev_status_w;
reg           csrbank17_ev_pending_re;
wire   [15:0] csrbank17_ev_pending_r;
reg           csrbank17_ev_pending_we;
wire   [15:0] csrbank17_ev_pending_w;
reg           csrbank17_ev_enable0_re;
wire   [15:0] csrbank17_ev_enable0_r;
reg           csrbank17_ev_enable0_we;
wire   [15:0] csrbank17_ev_enable0_w;
wire          csrbank17_sel;
wire          csrbank17_re;
wire   [15:0] interface18_bank_bus_adr;
wire          interface18_bank_bus_we;
wire   [31:0] interface18_bank_bus_dat_w;
reg    [31:0] interface18_bank_bus_dat_r;
wire          interface18_bank_bus_re;
reg           csrbank18_ev_soft0_re;
wire   [15:0] csrbank18_ev_soft0_r;
reg           csrbank18_ev_soft0_we;
wire   [15:0] csrbank18_ev_soft0_w;
reg           csrbank18_ev_edge_triggered0_re;
wire   [15:0] csrbank18_ev_edge_triggered0_r;
reg           csrbank18_ev_edge_triggered0_we;
wire   [15:0] csrbank18_ev_edge_triggered0_w;
reg           csrbank18_ev_polarity0_re;
wire   [15:0] csrbank18_ev_polarity0_r;
reg           csrbank18_ev_polarity0_we;
wire   [15:0] csrbank18_ev_polarity0_w;
reg           csrbank18_ev_status_re;
wire   [15:0] csrbank18_ev_status_r;
reg           csrbank18_ev_status_we;
wire   [15:0] csrbank18_ev_status_w;
reg           csrbank18_ev_pending_re;
wire   [15:0] csrbank18_ev_pending_r;
reg           csrbank18_ev_pending_we;
wire   [15:0] csrbank18_ev_pending_w;
reg           csrbank18_ev_enable0_re;
wire   [15:0] csrbank18_ev_enable0_r;
reg           csrbank18_ev_enable0_we;
wire   [15:0] csrbank18_ev_enable0_w;
wire          csrbank18_sel;
wire          csrbank18_re;
wire   [15:0] interface19_bank_bus_adr;
wire          interface19_bank_bus_we;
wire   [31:0] interface19_bank_bus_dat_w;
reg    [31:0] interface19_bank_bus_dat_r;
wire          interface19_bank_bus_re;
reg           csrbank19_ev_soft0_re;
wire   [15:0] csrbank19_ev_soft0_r;
reg           csrbank19_ev_soft0_we;
wire   [15:0] csrbank19_ev_soft0_w;
reg           csrbank19_ev_edge_triggered0_re;
wire   [15:0] csrbank19_ev_edge_triggered0_r;
reg           csrbank19_ev_edge_triggered0_we;
wire   [15:0] csrbank19_ev_edge_triggered0_w;
reg           csrbank19_ev_polarity0_re;
wire   [15:0] csrbank19_ev_polarity0_r;
reg           csrbank19_ev_polarity0_we;
wire   [15:0] csrbank19_ev_polarity0_w;
reg           csrbank19_ev_status_re;
wire   [15:0] csrbank19_ev_status_r;
reg           csrbank19_ev_status_we;
wire   [15:0] csrbank19_ev_status_w;
reg           csrbank19_ev_pending_re;
wire   [15:0] csrbank19_ev_pending_r;
reg           csrbank19_ev_pending_we;
wire   [15:0] csrbank19_ev_pending_w;
reg           csrbank19_ev_enable0_re;
wire   [15:0] csrbank19_ev_enable0_r;
reg           csrbank19_ev_enable0_we;
wire   [15:0] csrbank19_ev_enable0_w;
wire          csrbank19_sel;
wire          csrbank19_re;
wire   [15:0] interface20_bank_bus_adr;
wire          interface20_bank_bus_we;
wire   [31:0] interface20_bank_bus_dat_w;
reg    [31:0] interface20_bank_bus_dat_r;
wire          interface20_bank_bus_re;
reg           csrbank20_ev_soft0_re;
wire   [15:0] csrbank20_ev_soft0_r;
reg           csrbank20_ev_soft0_we;
wire   [15:0] csrbank20_ev_soft0_w;
reg           csrbank20_ev_edge_triggered0_re;
wire   [15:0] csrbank20_ev_edge_triggered0_r;
reg           csrbank20_ev_edge_triggered0_we;
wire   [15:0] csrbank20_ev_edge_triggered0_w;
reg           csrbank20_ev_polarity0_re;
wire   [15:0] csrbank20_ev_polarity0_r;
reg           csrbank20_ev_polarity0_we;
wire   [15:0] csrbank20_ev_polarity0_w;
reg           csrbank20_ev_status_re;
wire   [15:0] csrbank20_ev_status_r;
reg           csrbank20_ev_status_we;
wire   [15:0] csrbank20_ev_status_w;
reg           csrbank20_ev_pending_re;
wire   [15:0] csrbank20_ev_pending_r;
reg           csrbank20_ev_pending_we;
wire   [15:0] csrbank20_ev_pending_w;
reg           csrbank20_ev_enable0_re;
wire   [15:0] csrbank20_ev_enable0_r;
reg           csrbank20_ev_enable0_we;
wire   [15:0] csrbank20_ev_enable0_w;
wire          csrbank20_sel;
wire          csrbank20_re;
wire   [15:0] interface21_bank_bus_adr;
wire          interface21_bank_bus_we;
wire   [31:0] interface21_bank_bus_dat_w;
reg    [31:0] interface21_bank_bus_dat_r;
wire          interface21_bank_bus_re;
reg           csrbank21_ev_soft0_re;
wire   [15:0] csrbank21_ev_soft0_r;
reg           csrbank21_ev_soft0_we;
wire   [15:0] csrbank21_ev_soft0_w;
reg           csrbank21_ev_edge_triggered0_re;
wire   [15:0] csrbank21_ev_edge_triggered0_r;
reg           csrbank21_ev_edge_triggered0_we;
wire   [15:0] csrbank21_ev_edge_triggered0_w;
reg           csrbank21_ev_polarity0_re;
wire   [15:0] csrbank21_ev_polarity0_r;
reg           csrbank21_ev_polarity0_we;
wire   [15:0] csrbank21_ev_polarity0_w;
reg           csrbank21_ev_status_re;
wire   [15:0] csrbank21_ev_status_r;
reg           csrbank21_ev_status_we;
wire   [15:0] csrbank21_ev_status_w;
reg           csrbank21_ev_pending_re;
wire   [15:0] csrbank21_ev_pending_r;
reg           csrbank21_ev_pending_we;
wire   [15:0] csrbank21_ev_pending_w;
reg           csrbank21_ev_enable0_re;
wire   [15:0] csrbank21_ev_enable0_r;
reg           csrbank21_ev_enable0_we;
wire   [15:0] csrbank21_ev_enable0_w;
wire          csrbank21_sel;
wire          csrbank21_re;
wire   [15:0] interface22_bank_bus_adr;
wire          interface22_bank_bus_we;
wire   [31:0] interface22_bank_bus_dat_w;
reg    [31:0] interface22_bank_bus_dat_r;
wire          interface22_bank_bus_re;
reg           csrbank22_ev_soft0_re;
wire   [15:0] csrbank22_ev_soft0_r;
reg           csrbank22_ev_soft0_we;
wire   [15:0] csrbank22_ev_soft0_w;
reg           csrbank22_ev_edge_triggered0_re;
wire   [15:0] csrbank22_ev_edge_triggered0_r;
reg           csrbank22_ev_edge_triggered0_we;
wire   [15:0] csrbank22_ev_edge_triggered0_w;
reg           csrbank22_ev_polarity0_re;
wire   [15:0] csrbank22_ev_polarity0_r;
reg           csrbank22_ev_polarity0_we;
wire   [15:0] csrbank22_ev_polarity0_w;
reg           csrbank22_ev_status_re;
wire   [15:0] csrbank22_ev_status_r;
reg           csrbank22_ev_status_we;
wire   [15:0] csrbank22_ev_status_w;
reg           csrbank22_ev_pending_re;
wire   [15:0] csrbank22_ev_pending_r;
reg           csrbank22_ev_pending_we;
wire   [15:0] csrbank22_ev_pending_w;
reg           csrbank22_ev_enable0_re;
wire   [15:0] csrbank22_ev_enable0_r;
reg           csrbank22_ev_enable0_we;
wire   [15:0] csrbank22_ev_enable0_w;
wire          csrbank22_sel;
wire          csrbank22_re;
wire   [15:0] interface23_bank_bus_adr;
wire          interface23_bank_bus_we;
wire   [31:0] interface23_bank_bus_dat_w;
reg    [31:0] interface23_bank_bus_dat_r;
wire          interface23_bank_bus_re;
reg           csrbank23_wdata0_re;
wire   [31:0] csrbank23_wdata0_r;
reg           csrbank23_wdata0_we;
wire   [31:0] csrbank23_wdata0_w;
reg           csrbank23_rdata_re;
wire   [31:0] csrbank23_rdata_r;
reg           csrbank23_rdata_we;
wire   [31:0] csrbank23_rdata_w;
reg           csrbank23_ev_status_re;
wire    [3:0] csrbank23_ev_status_r;
reg           csrbank23_ev_status_we;
wire    [3:0] csrbank23_ev_status_w;
reg           csrbank23_ev_pending_re;
wire    [3:0] csrbank23_ev_pending_r;
reg           csrbank23_ev_pending_we;
wire    [3:0] csrbank23_ev_pending_w;
reg           csrbank23_ev_enable0_re;
wire    [3:0] csrbank23_ev_enable0_r;
reg           csrbank23_ev_enable0_we;
wire    [3:0] csrbank23_ev_enable0_w;
reg           csrbank23_status_re;
wire   [25:0] csrbank23_status_r;
reg           csrbank23_status_we;
wire   [25:0] csrbank23_status_w;
reg           csrbank23_control0_re;
wire          csrbank23_control0_r;
reg           csrbank23_control0_we;
wire          csrbank23_control0_w;
reg           csrbank23_done0_re;
wire          csrbank23_done0_r;
reg           csrbank23_done0_we;
wire          csrbank23_done0_w;
reg           csrbank23_loopback0_re;
wire          csrbank23_loopback0_r;
reg           csrbank23_loopback0_we;
wire          csrbank23_loopback0_w;
wire          csrbank23_sel;
wire          csrbank23_re;
wire   [15:0] interface24_bank_bus_adr;
wire          interface24_bank_bus_we;
wire   [31:0] interface24_bank_bus_dat_w;
reg    [31:0] interface24_bank_bus_dat_r;
wire          interface24_bank_bus_re;
reg           csrbank24_wdata0_re;
wire   [31:0] csrbank24_wdata0_r;
reg           csrbank24_wdata0_we;
wire   [31:0] csrbank24_wdata0_w;
reg           csrbank24_rdata_re;
wire   [31:0] csrbank24_rdata_r;
reg           csrbank24_rdata_we;
wire   [31:0] csrbank24_rdata_w;
reg           csrbank24_status_re;
wire    [5:0] csrbank24_status_r;
reg           csrbank24_status_we;
wire    [5:0] csrbank24_status_w;
reg           csrbank24_ev_status_re;
wire    [3:0] csrbank24_ev_status_r;
reg           csrbank24_ev_status_we;
wire    [3:0] csrbank24_ev_status_w;
reg           csrbank24_ev_pending_re;
wire    [3:0] csrbank24_ev_pending_r;
reg           csrbank24_ev_pending_we;
wire    [3:0] csrbank24_ev_pending_w;
reg           csrbank24_ev_enable0_re;
wire    [3:0] csrbank24_ev_enable0_r;
reg           csrbank24_ev_enable0_we;
wire    [3:0] csrbank24_ev_enable0_w;
reg           csrbank24_control0_re;
wire          csrbank24_control0_r;
reg           csrbank24_control0_we;
wire          csrbank24_control0_w;
reg           csrbank24_done0_re;
wire          csrbank24_done0_r;
reg           csrbank24_done0_we;
wire          csrbank24_done0_w;
wire          csrbank24_sel;
wire          csrbank24_re;
wire   [15:0] interface25_bank_bus_adr;
wire          interface25_bank_bus_we;
wire   [31:0] interface25_bank_bus_dat_w;
reg    [31:0] interface25_bank_bus_dat_r;
wire          interface25_bank_bus_re;
reg           csrbank25_pc_re;
wire   [31:0] csrbank25_pc_r;
reg           csrbank25_pc_we;
wire   [31:0] csrbank25_pc_w;
wire          csrbank25_sel;
wire          csrbank25_re;
wire   [15:0] interface26_bank_bus_adr;
wire          interface26_bank_bus_we;
wire   [31:0] interface26_bank_bus_dat_w;
reg    [31:0] interface26_bank_bus_dat_r;
wire          interface26_bank_bus_re;
reg           csrbank26_control0_re;
wire    [1:0] csrbank26_control0_r;
reg           csrbank26_control0_we;
wire    [1:0] csrbank26_control0_w;
reg           csrbank26_resume_time1_re;
wire   [31:0] csrbank26_resume_time1_r;
reg           csrbank26_resume_time1_we;
wire   [31:0] csrbank26_resume_time1_w;
reg           csrbank26_resume_time0_re;
wire   [31:0] csrbank26_resume_time0_r;
reg           csrbank26_resume_time0_we;
wire   [31:0] csrbank26_resume_time0_w;
reg           csrbank26_time1_re;
wire   [31:0] csrbank26_time1_r;
reg           csrbank26_time1_we;
wire   [31:0] csrbank26_time1_w;
reg           csrbank26_time0_re;
wire   [31:0] csrbank26_time0_r;
reg           csrbank26_time0_we;
wire   [31:0] csrbank26_time0_w;
reg           csrbank26_status_re;
wire          csrbank26_status_r;
reg           csrbank26_status_we;
wire          csrbank26_status_w;
reg           csrbank26_state0_re;
wire    [1:0] csrbank26_state0_r;
reg           csrbank26_state0_we;
wire    [1:0] csrbank26_state0_w;
reg           csrbank26_interrupt0_re;
wire          csrbank26_interrupt0_r;
reg           csrbank26_interrupt0_we;
wire          csrbank26_interrupt0_w;
reg           csrbank26_ev_status_re;
wire          csrbank26_ev_status_r;
reg           csrbank26_ev_status_we;
wire          csrbank26_ev_status_w;
reg           csrbank26_ev_pending_re;
wire          csrbank26_ev_pending_r;
reg           csrbank26_ev_pending_we;
wire          csrbank26_ev_pending_w;
reg           csrbank26_ev_enable0_re;
wire          csrbank26_ev_enable0_r;
reg           csrbank26_ev_enable0_we;
wire          csrbank26_ev_enable0_w;
wire          csrbank26_sel;
wire          csrbank26_re;
wire   [15:0] interface27_bank_bus_adr;
wire          interface27_bank_bus_we;
wire   [31:0] interface27_bank_bus_dat_w;
reg    [31:0] interface27_bank_bus_dat_r;
wire          interface27_bank_bus_re;
reg           csrbank27_control0_re;
wire          csrbank27_control0_r;
reg           csrbank27_control0_we;
wire          csrbank27_control0_w;
reg           csrbank27_time1_re;
wire   [31:0] csrbank27_time1_r;
reg           csrbank27_time1_we;
wire   [31:0] csrbank27_time1_w;
reg           csrbank27_time0_re;
wire   [31:0] csrbank27_time0_r;
reg           csrbank27_time0_we;
wire   [31:0] csrbank27_time0_w;
reg           csrbank27_msleep_target1_re;
wire   [31:0] csrbank27_msleep_target1_r;
reg           csrbank27_msleep_target1_we;
wire   [31:0] csrbank27_msleep_target1_w;
reg           csrbank27_msleep_target0_re;
wire   [31:0] csrbank27_msleep_target0_r;
reg           csrbank27_msleep_target0_we;
wire   [31:0] csrbank27_msleep_target0_w;
reg           csrbank27_ev_status_re;
wire          csrbank27_ev_status_r;
reg           csrbank27_ev_status_we;
wire          csrbank27_ev_status_w;
reg           csrbank27_ev_pending_re;
wire          csrbank27_ev_pending_r;
reg           csrbank27_ev_pending_we;
wire          csrbank27_ev_pending_w;
reg           csrbank27_ev_enable0_re;
wire          csrbank27_ev_enable0_r;
reg           csrbank27_ev_enable0_we;
wire          csrbank27_ev_enable0_w;
reg           csrbank27_clocks_per_tick0_re;
wire   [31:0] csrbank27_clocks_per_tick0_r;
reg           csrbank27_clocks_per_tick0_we;
wire   [31:0] csrbank27_clocks_per_tick0_w;
wire          csrbank27_sel;
wire          csrbank27_re;
wire   [15:0] interface28_bank_bus_adr;
wire          interface28_bank_bus_we;
wire   [31:0] interface28_bank_bus_dat_w;
reg    [31:0] interface28_bank_bus_dat_r;
wire          interface28_bank_bus_re;
reg           csrbank28_load0_re;
wire   [31:0] csrbank28_load0_r;
reg           csrbank28_load0_we;
wire   [31:0] csrbank28_load0_w;
reg           csrbank28_reload0_re;
wire   [31:0] csrbank28_reload0_r;
reg           csrbank28_reload0_we;
wire   [31:0] csrbank28_reload0_w;
reg           csrbank28_en0_re;
wire          csrbank28_en0_r;
reg           csrbank28_en0_we;
wire          csrbank28_en0_w;
reg           csrbank28_update_value0_re;
wire          csrbank28_update_value0_r;
reg           csrbank28_update_value0_we;
wire          csrbank28_update_value0_w;
reg           csrbank28_value_re;
wire   [31:0] csrbank28_value_r;
reg           csrbank28_value_we;
wire   [31:0] csrbank28_value_w;
reg           csrbank28_ev_status_re;
wire          csrbank28_ev_status_r;
reg           csrbank28_ev_status_we;
wire          csrbank28_ev_status_w;
reg           csrbank28_ev_pending_re;
wire          csrbank28_ev_pending_r;
reg           csrbank28_ev_pending_we;
wire          csrbank28_ev_pending_w;
reg           csrbank28_ev_enable0_re;
wire          csrbank28_ev_enable0_r;
reg           csrbank28_ev_enable0_we;
wire          csrbank28_ev_enable0_w;
wire          csrbank28_sel;
wire          csrbank28_re;
wire   [15:0] csr_interconnect_adr;
wire          csr_interconnect_we;
wire   [31:0] csr_interconnect_dat_w;
wire   [31:0] csr_interconnect_dat_r;
wire          csr_interconnect_re;
reg     [1:0] cramsoc_mailbox_state;
reg     [1:0] cramsoc_mailbox_next_state;
reg           mailbox_abort_ack1_mailbox_next_value0;
reg           mailbox_abort_ack1_mailbox_next_value_ce0;
reg           mailbox_abort_in_progress1_mailbox_next_value1;
reg           mailbox_abort_in_progress1_mailbox_next_value_ce1;
reg           mailbox_w_abort_mailbox_next_value2;
reg           mailbox_w_abort_mailbox_next_value_ce2;
reg     [1:0] cramsoc_mailboxclient_state;
reg     [1:0] cramsoc_mailboxclient_next_state;
reg           mb_client_abort_ack1_mailboxclient_next_value0;
reg           mb_client_abort_ack1_mailboxclient_next_value_ce0;
reg           mb_client_abort_in_progress1_mailboxclient_next_value1;
reg           mb_client_abort_in_progress1_mailboxclient_next_value_ce1;
reg           mb_client_w_abort_mailboxclient_next_value2;
reg           mb_client_w_abort_mailboxclient_next_value_ce2;
reg     [1:0] cramsoc_axilite2csr_state;
reg     [1:0] cramsoc_axilite2csr_next_state;
reg           cramsoc_last_was_read_axilite2csr_next_value;
reg           cramsoc_last_was_read_axilite2csr_next_value_ce;
wire   [29:0] slice_proxy0;
wire   [29:0] slice_proxy1;
reg           array_muxed0;
reg           array_muxed1;
reg           array_muxed2;
reg    [31:0] array_muxed3;
reg     [2:0] array_muxed4;
reg           array_muxed5;
reg           array_muxed6;
reg           array_muxed7;
reg    [31:0] array_muxed8;
reg     [3:0] array_muxed9;
reg           array_muxed10;
reg           array_muxed11;
reg           array_muxed12;
reg           array_muxed13;
reg    [31:0] array_muxed14;
reg     [2:0] array_muxed15;
reg           array_muxed16;
reg           multiregimpl0_regs0;
reg           multiregimpl0_regs1;
reg           multiregimpl1_regs0;
reg           multiregimpl1_regs1;
reg           multiregimpl2_regs0;
reg           multiregimpl2_regs1;
reg           multiregimpl3_regs0;
reg           multiregimpl3_regs1;
reg           multiregimpl4_regs0;
reg           multiregimpl4_regs1;
reg           multiregimpl5_regs0;
reg           multiregimpl5_regs1;
reg    [63:0] multiregimpl6_regs0;
reg    [63:0] multiregimpl6_regs1;
reg           multiregimpl7_regs0;
reg           multiregimpl7_regs1;
reg           multiregimpl8_regs0;
reg           multiregimpl8_regs1;
reg    [63:0] multiregimpl9_regs0;
reg    [63:0] multiregimpl9_regs1;
reg           multiregimpl10_regs0;
reg           multiregimpl10_regs1;
reg           multiregimpl11_regs0;
reg           multiregimpl11_regs1;
reg           multiregimpl12_regs0;
reg           multiregimpl12_regs1;
reg           multiregimpl13_regs0;
reg           multiregimpl13_regs1;
reg           multiregimpl14_regs0;
reg           multiregimpl14_regs1;
reg           multiregimpl15_regs0;
reg           multiregimpl15_regs1;
reg           multiregimpl16_regs0;
reg           multiregimpl16_regs1;
reg           multiregimpl17_regs0;
reg           multiregimpl17_regs1;
reg    [63:0] multiregimpl18_regs0;
reg    [63:0] multiregimpl18_regs1;

//------------------------------------------------------------------------------
// Combinatorial Logic
//------------------------------------------------------------------------------

assign sys_clk = aclk;
assign sys_rst = rst;
assign always_on_clk = always_on;
assign always_on_rst = sys_rst;
assign trimming_reset_1 = trimming_reset;
assign trimming_reset_ena_1 = trimming_reset_ena;
assign cramsoc_trimming_reset = trimming_reset_1;
assign cramsoc_trimming_reset_ena = trimming_reset_ena_1;
assign ibus_axi_awvalid = cramsoc_ibus_axi_aw_valid;
assign ibus_axi_awaddr = cramsoc_ibus_axi_aw_payload_addr;
assign ibus_axi_awburst = cramsoc_ibus_axi_aw_payload_burst;
assign ibus_axi_awlen = cramsoc_ibus_axi_aw_payload_len;
assign ibus_axi_awsize = cramsoc_ibus_axi_aw_payload_size;
assign ibus_axi_awlock = cramsoc_ibus_axi_aw_payload_lock;
assign ibus_axi_awprot = cramsoc_ibus_axi_aw_payload_prot;
assign ibus_axi_awcache = cramsoc_ibus_axi_aw_payload_cache;
assign ibus_axi_awqos = cramsoc_ibus_axi_aw_payload_qos;
assign ibus_axi_awregion = cramsoc_ibus_axi_aw_payload_region;
assign ibus_axi_awid = cramsoc_ibus_axi_aw_param_id;
assign ibus_axi_awuser = cramsoc_ibus_axi_aw_param_user;
assign cramsoc_ibus_axi_aw_ready = ibus_axi_awready;
assign ibus_axi_wvalid = cramsoc_ibus_axi_w_valid;
assign ibus_axi_wdata = cramsoc_ibus_axi_w_payload_data;
assign ibus_axi_wstrb = cramsoc_ibus_axi_w_payload_strb;
assign ibus_axi_wuser = cramsoc_ibus_axi_w_param_user;
assign ibus_axi_wlast = cramsoc_ibus_axi_w_last;
assign cramsoc_ibus_axi_w_ready = ibus_axi_wready;
assign cramsoc_ibus_axi_b_valid = ibus_axi_bvalid;
assign cramsoc_ibus_axi_b_payload_resp = ibus_axi_bresp;
assign cramsoc_ibus_axi_b_param_id = ibus_axi_bid;
assign cramsoc_ibus_axi_b_param_user = ibus_axi_buser;
assign ibus_axi_bready = cramsoc_ibus_axi_b_ready;
assign ibus_axi_arvalid = cramsoc_ibus_axi_ar_valid;
assign ibus_axi_araddr = cramsoc_ibus_axi_ar_payload_addr;
assign ibus_axi_arburst = cramsoc_ibus_axi_ar_payload_burst;
assign ibus_axi_arlen = cramsoc_ibus_axi_ar_payload_len;
assign ibus_axi_arsize = cramsoc_ibus_axi_ar_payload_size;
assign ibus_axi_arlock = cramsoc_ibus_axi_ar_payload_lock;
assign ibus_axi_arprot = cramsoc_ibus_axi_ar_payload_prot;
assign ibus_axi_arcache = cramsoc_ibus_axi_ar_payload_cache;
assign ibus_axi_arqos = cramsoc_ibus_axi_ar_payload_qos;
assign ibus_axi_arregion = cramsoc_ibus_axi_ar_payload_region;
assign ibus_axi_arid = cramsoc_ibus_axi_ar_param_id;
assign ibus_axi_aruser = cramsoc_ibus_axi_ar_param_user;
assign cramsoc_ibus_axi_ar_ready = ibus_axi_arready;
assign cramsoc_ibus_axi_r_valid = ibus_axi_rvalid;
assign cramsoc_ibus_axi_r_payload_resp = ibus_axi_rresp;
assign cramsoc_ibus_axi_r_payload_data = ibus_axi_rdata;
assign cramsoc_ibus_axi_r_param_id = ibus_axi_rid;
assign cramsoc_ibus_axi_r_param_user = ibus_axi_ruser;
assign cramsoc_ibus_axi_r_last = ibus_axi_rlast;
assign ibus_axi_rready = cramsoc_ibus_axi_r_ready;
assign dbus_axi_awvalid = cramsoc_dbus_aw_valid;
assign dbus_axi_awaddr = cramsoc_dbus_aw_payload_addr;
assign dbus_axi_awburst = cramsoc_dbus_aw_payload_burst;
assign dbus_axi_awlen = cramsoc_dbus_aw_payload_len;
assign dbus_axi_awsize = cramsoc_dbus_aw_payload_size;
assign dbus_axi_awlock = cramsoc_dbus_aw_payload_lock;
assign dbus_axi_awprot = cramsoc_dbus_aw_payload_prot;
assign dbus_axi_awcache = cramsoc_dbus_aw_payload_cache;
assign dbus_axi_awqos = cramsoc_dbus_aw_payload_qos;
assign dbus_axi_awregion = cramsoc_dbus_aw_payload_region;
assign dbus_axi_awid = cramsoc_dbus_aw_param_id;
assign dbus_axi_awuser = cramsoc_dbus_aw_param_user;
assign cramsoc_dbus_aw_ready = dbus_axi_awready;
assign dbus_axi_wvalid = cramsoc_dbus_w_valid;
assign dbus_axi_wdata = cramsoc_dbus_w_payload_data;
assign dbus_axi_wstrb = cramsoc_dbus_w_payload_strb;
assign dbus_axi_wuser = cramsoc_dbus_w_param_user;
assign dbus_axi_wlast = cramsoc_dbus_w_last;
assign cramsoc_dbus_w_ready = dbus_axi_wready;
assign cramsoc_dbus_b_valid = dbus_axi_bvalid;
assign cramsoc_dbus_b_payload_resp = dbus_axi_bresp;
assign cramsoc_dbus_b_param_id = dbus_axi_bid;
assign cramsoc_dbus_b_param_user = dbus_axi_buser;
assign dbus_axi_bready = cramsoc_dbus_b_ready;
assign dbus_axi_arvalid = cramsoc_dbus_ar_valid;
assign dbus_axi_araddr = cramsoc_dbus_ar_payload_addr;
assign dbus_axi_arburst = cramsoc_dbus_ar_payload_burst;
assign dbus_axi_arlen = cramsoc_dbus_ar_payload_len;
assign dbus_axi_arsize = cramsoc_dbus_ar_payload_size;
assign dbus_axi_arlock = cramsoc_dbus_ar_payload_lock;
assign dbus_axi_arprot = cramsoc_dbus_ar_payload_prot;
assign dbus_axi_arcache = cramsoc_dbus_ar_payload_cache;
assign dbus_axi_arqos = cramsoc_dbus_ar_payload_qos;
assign dbus_axi_arregion = cramsoc_dbus_ar_payload_region;
assign dbus_axi_arid = cramsoc_dbus_ar_param_id;
assign dbus_axi_aruser = cramsoc_dbus_ar_param_user;
assign cramsoc_dbus_ar_ready = dbus_axi_arready;
assign cramsoc_dbus_r_valid = dbus_axi_rvalid;
assign cramsoc_dbus_r_payload_resp = dbus_axi_rresp;
assign cramsoc_dbus_r_payload_data = dbus_axi_rdata;
assign cramsoc_dbus_r_param_id = dbus_axi_rid;
assign cramsoc_dbus_r_param_user = dbus_axi_ruser;
assign cramsoc_dbus_r_last = dbus_axi_rlast;
assign dbus_axi_rready = cramsoc_dbus_r_ready;
assign p_axi_awvalid = cramsoc_peripherals_aw_valid;
assign p_axi_awaddr = cramsoc_peripherals_aw_payload_addr;
assign p_axi_awprot = cramsoc_peripherals_aw_payload_prot;
assign cramsoc_peripherals_aw_ready = p_axi_awready;
assign p_axi_wvalid = cramsoc_peripherals_w_valid;
assign p_axi_wdata = cramsoc_peripherals_w_payload_data;
assign p_axi_wstrb = cramsoc_peripherals_w_payload_strb;
assign cramsoc_peripherals_w_ready = p_axi_wready;
assign cramsoc_peripherals_b_valid = p_axi_bvalid;
assign cramsoc_peripherals_b_payload_resp = p_axi_bresp;
assign p_axi_bready = cramsoc_peripherals_b_ready;
assign p_axi_arvalid = cramsoc_peripherals_ar_valid;
assign p_axi_araddr = cramsoc_peripherals_ar_payload_addr;
assign p_axi_arprot = cramsoc_peripherals_ar_payload_prot;
assign cramsoc_peripherals_ar_ready = p_axi_arready;
assign cramsoc_peripherals_r_valid = p_axi_rvalid;
assign cramsoc_peripherals_r_payload_resp = p_axi_rresp;
assign cramsoc_peripherals_r_payload_data = p_axi_rdata;
assign p_axi_rready = cramsoc_peripherals_r_ready;
assign cramsoc_cmbist = cmbist;
assign cramsoc_cmatpg = cmatpg;
assign cramsoc_vexsramtrm = vexsramtrm;
assign axi_active = ((((((((((((((((cramsoc_ibus_axi_ar_valid | cramsoc_ibus_axi_r_valid) | cramsoc_dbus_aw_valid) | cramsoc_dbus_w_valid) | cramsoc_dbus_b_valid) | cramsoc_dbus_ar_valid) | cramsoc_dbus_r_valid) | cramsoc_peripherals_aw_valid) | cramsoc_peripherals_w_valid) | cramsoc_peripherals_b_valid) | cramsoc_peripherals_ar_valid) | cramsoc_peripherals_r_valid) | ibus_r_active) | dbus_r_active) | dbus_w_active) | pbus_r_active) | pbus_w_active);
assign sleep_req = (((cramsoc_wfi_active & cpu_int_active) & (~axi_active)) & (active_timeout == 1'd0));
always @(*) begin
    irq_remap0 <= 16'd0;
    irq_remap0[0] <= irqarray_bank2[1];
    irq_remap0[1] <= irqarray_bank0[1];
    irq_remap0[2] <= irqarray_bank0[2];
    irq_remap0[3] <= irqarray_bank0[3];
    irq_remap0[4] <= irqarray_bank10[3];
    irq_remap0[5] <= irqarray_bank10[4];
    irq_remap0[6] <= irqarray_bank10[5];
    irq_remap0[7] <= irqarray_bank10[6];
    irq_remap0[8] <= irqarray_bank0[8];
    irq_remap0[9] <= irqarray_bank0[9];
    irq_remap0[10] <= irqarray_bank0[10];
    irq_remap0[11] <= irqarray_bank0[11];
    irq_remap0[12] <= irqarray_bank0[12];
    irq_remap0[13] <= irqarray_bank0[13];
    irq_remap0[14] <= irqarray_bank0[14];
    irq_remap0[15] <= irqarray_bank0[15];
end
always @(*) begin
    irq_remap1 <= 16'd0;
    irq_remap1[0] <= irqarray_bank10[1];
    irq_remap1[1] <= irqarray_bank1[1];
    irq_remap1[2] <= irqarray_bank1[2];
    irq_remap1[3] <= irqarray_bank1[3];
    irq_remap1[4] <= irqarray_bank1[4];
    irq_remap1[5] <= irqarray_bank1[5];
    irq_remap1[6] <= irqarray_bank1[6];
    irq_remap1[7] <= irqarray_bank1[7];
    irq_remap1[8] <= irqarray_bank1[8];
    irq_remap1[9] <= irqarray_bank1[9];
    irq_remap1[10] <= irqarray_bank1[10];
    irq_remap1[11] <= irqarray_bank1[11];
    irq_remap1[12] <= irqarray_bank1[12];
    irq_remap1[13] <= irqarray_bank1[13];
    irq_remap1[14] <= irqarray_bank1[14];
    irq_remap1[15] <= irqarray_bank1[15];
end
always @(*) begin
    irq_remap2 <= 16'd0;
    irq_remap2[0] <= irqarray_bank2[0];
    irq_remap2[1] <= irqarray_bank2[1];
    irq_remap2[2] <= irqarray_bank2[2];
    irq_remap2[3] <= irqarray_bank2[3];
    irq_remap2[4] <= irqarray_bank2[4];
    irq_remap2[5] <= irqarray_bank2[5];
    irq_remap2[6] <= irqarray_bank2[6];
    irq_remap2[7] <= irqarray_bank2[7];
    irq_remap2[8] <= irqarray_bank2[8];
    irq_remap2[9] <= irqarray_bank2[9];
    irq_remap2[10] <= irqarray_bank2[10];
    irq_remap2[11] <= irqarray_bank2[11];
    irq_remap2[12] <= irqarray_bank2[12];
    irq_remap2[13] <= irqarray_bank2[13];
    irq_remap2[14] <= irqarray_bank2[14];
    irq_remap2[15] <= irqarray_bank2[15];
end
always @(*) begin
    irq_remap3 <= 16'd0;
    irq_remap3[0] <= irqarray_bank3[0];
    irq_remap3[1] <= irqarray_bank3[1];
    irq_remap3[2] <= irqarray_bank3[2];
    irq_remap3[3] <= irqarray_bank3[3];
    irq_remap3[4] <= irqarray_bank3[4];
    irq_remap3[5] <= irqarray_bank3[5];
    irq_remap3[6] <= irqarray_bank3[6];
    irq_remap3[7] <= irqarray_bank3[7];
    irq_remap3[8] <= irqarray_bank3[8];
    irq_remap3[9] <= irqarray_bank3[9];
    irq_remap3[10] <= irqarray_bank3[10];
    irq_remap3[11] <= irqarray_bank3[11];
    irq_remap3[12] <= irqarray_bank3[12];
    irq_remap3[13] <= irqarray_bank3[13];
    irq_remap3[14] <= irqarray_bank3[14];
    irq_remap3[15] <= irqarray_bank3[15];
end
always @(*) begin
    irq_remap4 <= 16'd0;
    irq_remap4[0] <= irqarray_bank3[0];
    irq_remap4[1] <= irqarray_bank3[1];
    irq_remap4[2] <= irqarray_bank3[2];
    irq_remap4[3] <= irqarray_bank3[3];
    irq_remap4[4] <= irqarray_bank3[4];
    irq_remap4[5] <= irqarray_bank3[5];
    irq_remap4[6] <= irqarray_bank3[6];
    irq_remap4[7] <= irqarray_bank3[7];
    irq_remap4[8] <= irqarray_bank4[8];
    irq_remap4[9] <= irqarray_bank4[9];
    irq_remap4[10] <= irqarray_bank4[10];
    irq_remap4[11] <= irqarray_bank4[11];
    irq_remap4[12] <= irqarray_bank4[12];
    irq_remap4[13] <= irqarray_bank4[13];
    irq_remap4[14] <= irqarray_bank4[14];
    irq_remap4[15] <= irqarray_bank4[15];
end
always @(*) begin
    irq_remap5 <= 16'd0;
    irq_remap5[0] <= irqarray_bank5[0];
    irq_remap5[1] <= irqarray_bank5[1];
    irq_remap5[2] <= irqarray_bank5[2];
    irq_remap5[3] <= irqarray_bank5[3];
    irq_remap5[4] <= irqarray_bank5[4];
    irq_remap5[5] <= irqarray_bank5[5];
    irq_remap5[6] <= irqarray_bank5[6];
    irq_remap5[7] <= irqarray_bank5[7];
    irq_remap5[8] <= irqarray_bank5[8];
    irq_remap5[9] <= irqarray_bank5[9];
    irq_remap5[10] <= irqarray_bank5[10];
    irq_remap5[11] <= irqarray_bank5[11];
    irq_remap5[12] <= irqarray_bank5[12];
    irq_remap5[13] <= irqarray_bank5[13];
    irq_remap5[14] <= irqarray_bank5[14];
    irq_remap5[15] <= irqarray_bank5[15];
end
always @(*) begin
    irq_remap6 <= 16'd0;
    irq_remap6[0] <= irqarray_bank6[0];
    irq_remap6[1] <= irqarray_bank6[1];
    irq_remap6[2] <= irqarray_bank6[2];
    irq_remap6[3] <= irqarray_bank6[3];
    irq_remap6[4] <= irqarray_bank6[4];
    irq_remap6[5] <= irqarray_bank6[5];
    irq_remap6[6] <= irqarray_bank6[6];
    irq_remap6[7] <= irqarray_bank6[7];
    irq_remap6[8] <= irqarray_bank6[8];
    irq_remap6[9] <= irqarray_bank6[9];
    irq_remap6[10] <= irqarray_bank6[10];
    irq_remap6[11] <= irqarray_bank6[11];
    irq_remap6[12] <= irqarray_bank6[12];
    irq_remap6[13] <= irqarray_bank6[13];
    irq_remap6[14] <= irqarray_bank6[14];
    irq_remap6[15] <= irqarray_bank6[15];
end
always @(*) begin
    irq_remap7 <= 16'd0;
    irq_remap7[0] <= irqarray_bank7[0];
    irq_remap7[1] <= irqarray_bank7[1];
    irq_remap7[2] <= irqarray_bank7[2];
    irq_remap7[3] <= irqarray_bank7[3];
    irq_remap7[4] <= irqarray_bank7[4];
    irq_remap7[5] <= irqarray_bank7[5];
    irq_remap7[6] <= irqarray_bank7[6];
    irq_remap7[7] <= irqarray_bank7[7];
    irq_remap7[8] <= irqarray_bank7[8];
    irq_remap7[9] <= irqarray_bank7[9];
    irq_remap7[10] <= irqarray_bank7[10];
    irq_remap7[11] <= irqarray_bank7[11];
    irq_remap7[12] <= irqarray_bank7[12];
    irq_remap7[13] <= irqarray_bank7[13];
    irq_remap7[14] <= irqarray_bank7[14];
    irq_remap7[15] <= irqarray_bank7[15];
end
always @(*) begin
    irq_remap8 <= 16'd0;
    irq_remap8[0] <= irqarray_bank8[0];
    irq_remap8[1] <= irqarray_bank8[1];
    irq_remap8[2] <= irqarray_bank8[2];
    irq_remap8[3] <= irqarray_bank8[3];
    irq_remap8[4] <= irqarray_bank8[4];
    irq_remap8[5] <= irqarray_bank8[5];
    irq_remap8[6] <= irqarray_bank8[6];
    irq_remap8[7] <= irqarray_bank8[7];
    irq_remap8[8] <= irqarray_bank8[8];
    irq_remap8[9] <= irqarray_bank8[9];
    irq_remap8[10] <= irqarray_bank8[10];
    irq_remap8[11] <= irqarray_bank8[11];
    irq_remap8[12] <= irqarray_bank8[12];
    irq_remap8[13] <= irqarray_bank8[13];
    irq_remap8[14] <= irqarray_bank8[14];
    irq_remap8[15] <= irqarray_bank8[15];
end
always @(*) begin
    irq_remap9 <= 16'd0;
    irq_remap9[0] <= irqarray_bank9[0];
    irq_remap9[1] <= irqarray_bank9[1];
    irq_remap9[2] <= irqarray_bank9[2];
    irq_remap9[3] <= irqarray_bank9[3];
    irq_remap9[4] <= irqarray_bank9[4];
    irq_remap9[5] <= irqarray_bank9[5];
    irq_remap9[6] <= irqarray_bank9[6];
    irq_remap9[7] <= irqarray_bank9[7];
    irq_remap9[8] <= irqarray_bank9[8];
    irq_remap9[9] <= irqarray_bank9[9];
    irq_remap9[10] <= irqarray_bank9[10];
    irq_remap9[11] <= irqarray_bank9[11];
    irq_remap9[12] <= irqarray_bank9[12];
    irq_remap9[13] <= irqarray_bank9[13];
    irq_remap9[14] <= irqarray_bank9[14];
    irq_remap9[15] <= irqarray_bank9[15];
end
always @(*) begin
    irq_remap10 <= 16'd0;
    irq_remap10[0] <= irqarray_bank10[0];
    irq_remap10[1] <= irqarray_bank10[1];
    irq_remap10[2] <= irqarray_bank10[2];
    irq_remap10[3] <= irqarray_bank10[3];
    irq_remap10[4] <= irqarray_bank10[4];
    irq_remap10[5] <= irqarray_bank10[5];
    irq_remap10[6] <= irqarray_bank10[6];
    irq_remap10[7] <= irqarray_bank10[7];
    irq_remap10[8] <= irqarray_bank10[8];
    irq_remap10[9] <= irqarray_bank10[9];
    irq_remap10[10] <= irqarray_bank10[10];
    irq_remap10[11] <= irqarray_bank10[11];
    irq_remap10[12] <= irqarray_bank10[12];
    irq_remap10[13] <= irqarray_bank10[13];
    irq_remap10[14] <= irqarray_bank10[14];
    irq_remap10[15] <= irqarray_bank10[15];
end
always @(*) begin
    irq_remap11 <= 16'd0;
    irq_remap11[0] <= irqarray_bank8[4];
    irq_remap11[1] <= irqarray_bank8[5];
    irq_remap11[2] <= irqarray_bank11[2];
    irq_remap11[3] <= irqarray_bank11[3];
    irq_remap11[4] <= irqarray_bank11[4];
    irq_remap11[5] <= irqarray_bank11[5];
    irq_remap11[6] <= irqarray_bank11[6];
    irq_remap11[7] <= irqarray_bank11[7];
    irq_remap11[8] <= irqarray_bank11[8];
    irq_remap11[9] <= irqarray_bank11[9];
    irq_remap11[10] <= irqarray_bank11[10];
    irq_remap11[11] <= irqarray_bank11[11];
    irq_remap11[12] <= irqarray_bank11[12];
    irq_remap11[13] <= irqarray_bank11[13];
    irq_remap11[14] <= irqarray_bank11[14];
    irq_remap11[15] <= irqarray_bank11[15];
end
always @(*) begin
    irq_remap12 <= 16'd0;
    irq_remap12[0] <= irqarray_bank12[0];
    irq_remap12[1] <= irqarray_bank12[1];
    irq_remap12[2] <= irqarray_bank12[2];
    irq_remap12[3] <= irqarray_bank12[3];
    irq_remap12[4] <= irqarray_bank12[4];
    irq_remap12[5] <= irqarray_bank12[5];
    irq_remap12[6] <= irqarray_bank12[6];
    irq_remap12[7] <= irqarray_bank12[7];
    irq_remap12[8] <= irqarray_bank12[8];
    irq_remap12[9] <= irqarray_bank12[9];
    irq_remap12[10] <= irqarray_bank12[10];
    irq_remap12[11] <= irqarray_bank12[11];
    irq_remap12[12] <= irqarray_bank12[12];
    irq_remap12[13] <= irqarray_bank12[13];
    irq_remap12[14] <= irqarray_bank12[14];
    irq_remap12[15] <= irqarray_bank12[15];
end
always @(*) begin
    irq_remap13 <= 16'd0;
    irq_remap13[0] <= irqarray_bank13[0];
    irq_remap13[1] <= irqarray_bank13[1];
    irq_remap13[2] <= irqarray_bank13[2];
    irq_remap13[3] <= irqarray_bank13[3];
    irq_remap13[4] <= irqarray_bank13[4];
    irq_remap13[5] <= irqarray_bank13[5];
    irq_remap13[6] <= irqarray_bank13[6];
    irq_remap13[7] <= irqarray_bank13[7];
    irq_remap13[8] <= irqarray_bank13[8];
    irq_remap13[9] <= irqarray_bank13[9];
    irq_remap13[10] <= irqarray_bank13[10];
    irq_remap13[11] <= irqarray_bank13[11];
    irq_remap13[12] <= irqarray_bank13[12];
    irq_remap13[13] <= irqarray_bank13[13];
    irq_remap13[14] <= irqarray_bank13[14];
    irq_remap13[15] <= irqarray_bank13[15];
end
always @(*) begin
    irq_remap14 <= 16'd0;
    irq_remap14[0] <= irqarray_bank5[8];
    irq_remap14[1] <= irqarray_bank5[9];
    irq_remap14[2] <= irqarray_bank5[10];
    irq_remap14[3] <= irqarray_bank5[11];
    irq_remap14[4] <= irqarray_bank5[12];
    irq_remap14[5] <= irqarray_bank5[13];
    irq_remap14[6] <= irqarray_bank5[14];
    irq_remap14[7] <= irqarray_bank5[15];
    irq_remap14[8] <= irqarray_bank3[0];
    irq_remap14[9] <= irqarray_bank14[9];
    irq_remap14[10] <= irqarray_bank14[10];
    irq_remap14[11] <= irqarray_bank14[11];
    irq_remap14[12] <= irqarray_bank14[12];
    irq_remap14[13] <= irqarray_bank14[13];
    irq_remap14[14] <= irqarray_bank14[14];
    irq_remap14[15] <= irqarray_bank14[15];
end
always @(*) begin
    irq_remap15 <= 16'd0;
    irq_remap15[0] <= irqarray_bank15[0];
    irq_remap15[1] <= irqarray_bank15[1];
    irq_remap15[2] <= irqarray_bank15[2];
    irq_remap15[3] <= irqarray_bank15[3];
    irq_remap15[4] <= irqarray_bank15[4];
    irq_remap15[5] <= irqarray_bank15[5];
    irq_remap15[6] <= irqarray_bank15[6];
    irq_remap15[7] <= irqarray_bank15[7];
    irq_remap15[8] <= irqarray_bank15[8];
    irq_remap15[9] <= irqarray_bank15[9];
    irq_remap15[10] <= irqarray_bank15[10];
    irq_remap15[11] <= irqarray_bank15[11];
    irq_remap15[12] <= irqarray_bank15[12];
    irq_remap15[13] <= irqarray_bank15[13];
    irq_remap15[14] <= irqarray_bank15[14];
    irq_remap15[15] <= irqarray_bank15[15];
end
always @(*) begin
    irq_remap16 <= 16'd0;
    irq_remap16[0] <= irqarray_bank8[8];
    irq_remap16[1] <= irqarray_bank8[4];
    irq_remap16[2] <= irqarray_bank8[5];
    irq_remap16[3] <= irqarray_bank16[3];
    irq_remap16[4] <= irqarray_bank6[4];
    irq_remap16[5] <= irqarray_bank6[5];
    irq_remap16[6] <= irqarray_bank6[6];
    irq_remap16[7] <= irqarray_bank6[7];
    irq_remap16[8] <= irqarray_bank6[8];
    irq_remap16[9] <= irqarray_bank6[9];
    irq_remap16[10] <= irqarray_bank6[10];
    irq_remap16[11] <= irqarray_bank6[11];
    irq_remap16[12] <= irqarray_bank7[0];
    irq_remap16[13] <= irqarray_bank7[1];
    irq_remap16[14] <= irqarray_bank7[2];
    irq_remap16[15] <= irqarray_bank7[3];
end
always @(*) begin
    irq_remap17 <= 16'd0;
    irq_remap17[0] <= irqarray_bank7[4];
    irq_remap17[1] <= irqarray_bank7[5];
    irq_remap17[2] <= irqarray_bank7[6];
    irq_remap17[3] <= irqarray_bank7[7];
    irq_remap17[4] <= irqarray_bank10[3];
    irq_remap17[5] <= irqarray_bank10[4];
    irq_remap17[6] <= irqarray_bank10[5];
    irq_remap17[7] <= irqarray_bank10[6];
    irq_remap17[8] <= irqarray_bank2[0];
    irq_remap17[9] <= irqarray_bank8[9];
    irq_remap17[10] <= irqarray_bank10[0];
    irq_remap17[11] <= irqarray_bank10[2];
    irq_remap17[12] <= irqarray_bank17[12];
    irq_remap17[13] <= irqarray_bank17[13];
    irq_remap17[14] <= irqarray_bank17[14];
    irq_remap17[15] <= irqarray_bank17[15];
end
always @(*) begin
    irq_remap18 <= 16'd0;
    irq_remap18[0] <= irqarray_bank10[3];
    irq_remap18[1] <= irqarray_bank10[4];
    irq_remap18[2] <= irqarray_bank10[5];
    irq_remap18[3] <= irqarray_bank10[6];
    irq_remap18[4] <= irqarray_bank7[8];
    irq_remap18[5] <= irqarray_bank7[9];
    irq_remap18[6] <= irqarray_bank7[10];
    irq_remap18[7] <= irqarray_bank7[11];
    irq_remap18[8] <= irqarray_bank12[8];
    irq_remap18[9] <= irqarray_bank12[9];
    irq_remap18[10] <= irqarray_bank12[10];
    irq_remap18[11] <= irqarray_bank12[12];
    irq_remap18[12] <= irqarray_bank12[13];
    irq_remap18[13] <= irqarray_bank12[14];
    irq_remap18[14] <= irqarray_bank10[0];
    irq_remap18[15] <= irqarray_bank8[8];
end
always @(*) begin
    irq_remap19 <= 16'd0;
    irq_remap19[0] <= irqarray_bank2[2];
    irq_remap19[1] <= irqarray_bank2[3];
    irq_remap19[2] <= irqarray_bank2[4];
    irq_remap19[3] <= irqarray_bank2[5];
    irq_remap19[4] <= irqarray_bank10[3];
    irq_remap19[5] <= irqarray_bank10[4];
    irq_remap19[6] <= irqarray_bank10[5];
    irq_remap19[7] <= irqarray_bank10[6];
    irq_remap19[8] <= irqarray_bank8[0];
    irq_remap19[9] <= irqarray_bank8[1];
    irq_remap19[10] <= irqarray_bank8[2];
    irq_remap19[11] <= irqarray_bank8[3];
    irq_remap19[12] <= irqarray_bank19[12];
    irq_remap19[13] <= irqarray_bank19[13];
    irq_remap19[14] <= irqarray_bank19[14];
    irq_remap19[15] <= irqarray_bank19[15];
end
assign susres_time_status = ticktimer_timer1;
assign susres_paused = ticktimer_paused0;
assign ticktimer_resume_time = susres_resume_time_storage;
assign ticktimer_pause0 = susres_pause;
assign ticktimer_load = susres_load;
assign mailbox_cmatpg = cmatpg;
assign mailbox_cmbist = cmbist;
assign mailbox_vexsramtrm = vexsramtrm;
assign loopback = mailbox_loopback;
assign mailbox_reset_n = (~sys_rst);
assign w_dat = mailbox_w_dat;
assign w_valid = mailbox_w_valid;
assign w_done = mailbox_w_done;
assign mailbox_w_ready = w_ready;
assign mailbox_r_dat = r_dat;
assign mailbox_r_valid = r_valid;
assign mailbox_r_done = r_done;
assign r_ready = mailbox_r_ready;
assign mailbox_r_abort = r_abort;
assign w_abort = mailbox_w_abort;
always @(*) begin
    r_dat <= 32'd0;
    r_valid <= 1'd0;
    r_done <= 1'd0;
    mb_client_reset_n <= 1'd0;
    r_abort <= 1'd0;
    w_ready <= 1'd0;
    if (loopback) begin
        mb_client_reset_n <= (~sys_rst);
        r_dat <= mb_client_w_dat;
        r_valid <= mb_client_w_valid;
        r_done <= mb_client_w_done;
        w_ready <= mb_client_r_ready;
        r_abort <= mb_client_w_abort;
    end else begin
        r_dat <= mbox_w_dat;
        r_valid <= mbox_w_valid;
        r_done <= mbox_w_done;
        w_ready <= mbox_r_ready;
        r_abort <= mbox_w_abort;
    end
end
assign mb_client_w_ready = r_ready;
assign mb_client_r_dat = w_dat;
assign mb_client_r_valid = w_valid;
assign mb_client_r_done = w_done;
assign mb_client_r_abort = w_abort;
assign mbox_w_ready = r_ready;
assign mbox_r_dat = w_dat;
assign mbox_r_valid = w_valid;
assign mbox_r_done = w_done;
assign mbox_r_abort = w_abort;
assign test = csr_wtest_storage;
always @(*) begin
    cramsoc_interrupt <= 32'd0;
    cramsoc_interrupt[0] <= irqarray0_irq;
    cramsoc_interrupt[1] <= irqarray1_irq;
    cramsoc_interrupt[10] <= irqarray10_irq;
    cramsoc_interrupt[11] <= irqarray11_irq;
    cramsoc_interrupt[12] <= irqarray12_irq;
    cramsoc_interrupt[13] <= irqarray13_irq;
    cramsoc_interrupt[14] <= irqarray14_irq;
    cramsoc_interrupt[15] <= irqarray15_irq;
    cramsoc_interrupt[16] <= irqarray16_irq;
    cramsoc_interrupt[17] <= irqarray17_irq;
    cramsoc_interrupt[18] <= irqarray18_irq;
    cramsoc_interrupt[19] <= irqarray19_irq;
    cramsoc_interrupt[2] <= irqarray2_irq;
    cramsoc_interrupt[3] <= irqarray3_irq;
    cramsoc_interrupt[4] <= irqarray4_irq;
    cramsoc_interrupt[5] <= irqarray5_irq;
    cramsoc_interrupt[6] <= irqarray6_irq;
    cramsoc_interrupt[7] <= irqarray7_irq;
    cramsoc_interrupt[8] <= irqarray8_irq;
    cramsoc_interrupt[9] <= irqarray9_irq;
    cramsoc_interrupt[22] <= mailbox_irq;
    cramsoc_interrupt[23] <= mb_client_irq;
    cramsoc_interrupt[21] <= susres_irq;
    cramsoc_interrupt[20] <= ticktimer_irq;
    cramsoc_interrupt[30] <= cramsoc_irq;
end
assign socbushandler_slave_sel_dec0 = (slice_proxy0[29:16] == 14'd14336);
assign socbushandler_slave_sel_dec1 = (slice_proxy1[29:16] == 14'd14336);
always @(*) begin
    socbushandler_slave_sel0 <= 1'd0;
    if (socbushandler_axiliterequestcounter0_empty) begin
        socbushandler_slave_sel0 <= socbushandler_slave_sel_dec0;
    end else begin
        socbushandler_slave_sel0 <= socbushandler_slave_sel_reg0;
    end
end
always @(*) begin
    socbushandler_slave_sel1 <= 1'd0;
    if (socbushandler_axiliterequestcounter1_empty) begin
        socbushandler_slave_sel1 <= socbushandler_slave_sel_dec1;
    end else begin
        socbushandler_slave_sel1 <= socbushandler_slave_sel_reg1;
    end
end
assign socbushandler_aw_valid = (cramsoc_corecsr_aw_valid & socbushandler_slave_sel0);
assign socbushandler_aw_first = cramsoc_corecsr_aw_first;
assign socbushandler_aw_last = cramsoc_corecsr_aw_last;
assign socbushandler_aw_payload_addr = cramsoc_corecsr_aw_payload_addr;
assign socbushandler_aw_payload_prot = cramsoc_corecsr_aw_payload_prot;
assign socbushandler_w_valid = (cramsoc_corecsr_w_valid & socbushandler_slave_sel0);
assign socbushandler_w_first = cramsoc_corecsr_w_first;
assign socbushandler_w_last = cramsoc_corecsr_w_last;
assign socbushandler_w_payload_data = cramsoc_corecsr_w_payload_data;
assign socbushandler_w_payload_strb = cramsoc_corecsr_w_payload_strb;
assign socbushandler_b_ready = (cramsoc_corecsr_b_ready & socbushandler_slave_sel0);
assign socbushandler_ar_valid = (cramsoc_corecsr_ar_valid & socbushandler_slave_sel1);
assign socbushandler_ar_first = cramsoc_corecsr_ar_first;
assign socbushandler_ar_last = cramsoc_corecsr_ar_last;
assign socbushandler_ar_payload_addr = cramsoc_corecsr_ar_payload_addr;
assign socbushandler_ar_payload_prot = cramsoc_corecsr_ar_payload_prot;
assign socbushandler_r_ready = (cramsoc_corecsr_r_ready & socbushandler_slave_sel1);
assign cramsoc_corecsr_aw_ready = (socbushandler_aw_ready & {1{socbushandler_slave_sel0}});
assign cramsoc_corecsr_w_ready = (socbushandler_w_ready & {1{socbushandler_slave_sel0}});
assign cramsoc_corecsr_b_valid = (socbushandler_b_valid & {1{socbushandler_slave_sel0}});
assign cramsoc_corecsr_b_first = (socbushandler_b_first & {1{socbushandler_slave_sel0}});
assign cramsoc_corecsr_b_last = (socbushandler_b_last & {1{socbushandler_slave_sel0}});
assign cramsoc_corecsr_b_payload_resp = (socbushandler_b_payload_resp & {2{socbushandler_slave_sel0}});
assign cramsoc_corecsr_ar_ready = (socbushandler_ar_ready & {1{socbushandler_slave_sel1}});
assign cramsoc_corecsr_r_valid = (socbushandler_r_valid & {1{socbushandler_slave_sel1}});
assign cramsoc_corecsr_r_first = (socbushandler_r_first & {1{socbushandler_slave_sel1}});
assign cramsoc_corecsr_r_last = (socbushandler_r_last & {1{socbushandler_slave_sel1}});
assign cramsoc_corecsr_r_payload_resp = (socbushandler_r_payload_resp & {2{socbushandler_slave_sel1}});
assign cramsoc_corecsr_r_payload_data = (socbushandler_r_payload_data & {32{socbushandler_slave_sel1}});
assign socbushandler_axiliterequestcounter0_full = (socbushandler_axiliterequestcounter0_counter == 8'd255);
assign socbushandler_axiliterequestcounter0_empty = (socbushandler_axiliterequestcounter0_counter == 1'd0);
assign socbushandler_axiliterequestcounter0_stall = ((cramsoc_corecsr_aw_valid & cramsoc_corecsr_aw_ready) & socbushandler_axiliterequestcounter0_full);
assign socbushandler_axiliterequestcounter1_full = (socbushandler_axiliterequestcounter1_counter == 8'd255);
assign socbushandler_axiliterequestcounter1_empty = (socbushandler_axiliterequestcounter1_counter == 1'd0);
assign socbushandler_axiliterequestcounter1_stall = ((cramsoc_corecsr_ar_valid & cramsoc_corecsr_ar_ready) & socbushandler_axiliterequestcounter1_full);
assign cramsoc_aw_valid = array_muxed0;
assign cramsoc_aw_first = array_muxed1;
assign cramsoc_aw_last = array_muxed2;
assign cramsoc_aw_payload_addr = array_muxed3;
assign cramsoc_aw_payload_prot = array_muxed4;
assign cramsoc_w_valid = array_muxed5;
assign cramsoc_w_first = array_muxed6;
assign cramsoc_w_last = array_muxed7;
assign cramsoc_w_payload_data = array_muxed8;
assign cramsoc_w_payload_strb = array_muxed9;
assign cramsoc_b_ready = array_muxed10;
assign cramsoc_ar_valid = array_muxed11;
assign cramsoc_ar_first = array_muxed12;
assign cramsoc_ar_last = array_muxed13;
assign cramsoc_ar_payload_addr = array_muxed14;
assign cramsoc_ar_payload_prot = array_muxed15;
assign cramsoc_r_ready = array_muxed16;
always @(*) begin
    socbushandler_aw_ready <= 1'd0;
    if ((socbushandler_rr_write_grant == 1'd0)) begin
        socbushandler_aw_ready <= cramsoc_aw_ready;
    end
end
always @(*) begin
    socbushandler_w_ready <= 1'd0;
    if ((socbushandler_rr_write_grant == 1'd0)) begin
        socbushandler_w_ready <= cramsoc_w_ready;
    end
end
always @(*) begin
    socbushandler_b_valid <= 1'd0;
    if ((socbushandler_rr_write_grant == 1'd0)) begin
        socbushandler_b_valid <= cramsoc_b_valid;
    end
end
assign socbushandler_b_first = cramsoc_b_first;
assign socbushandler_b_last = cramsoc_b_last;
assign socbushandler_b_payload_resp = cramsoc_b_payload_resp;
always @(*) begin
    socbushandler_ar_ready <= 1'd0;
    if ((socbushandler_rr_read_grant == 1'd0)) begin
        socbushandler_ar_ready <= cramsoc_ar_ready;
    end
end
always @(*) begin
    socbushandler_r_valid <= 1'd0;
    if ((socbushandler_rr_read_grant == 1'd0)) begin
        socbushandler_r_valid <= cramsoc_r_valid;
    end
end
assign socbushandler_r_first = cramsoc_r_first;
assign socbushandler_r_last = cramsoc_r_last;
assign socbushandler_r_payload_resp = cramsoc_r_payload_resp;
assign socbushandler_r_payload_data = cramsoc_r_payload_data;
assign socbushandler_rr_write_ce = ((~((cramsoc_aw_valid | cramsoc_w_valid) | cramsoc_b_valid)) & socbushandler_wr_lock_empty);
assign socbushandler_rr_read_ce = ((~(cramsoc_ar_valid | cramsoc_r_valid)) & socbushandler_rd_lock_empty);
assign socbushandler_rr_write_request = {((socbushandler_aw_valid | socbushandler_w_valid) | socbushandler_b_valid)};
assign socbushandler_rr_read_request = {(socbushandler_ar_valid | socbushandler_r_valid)};
assign socbushandler_rr_write_grant = 1'd0;
assign socbushandler_rr_read_grant = 1'd0;
assign socbushandler_wr_lock_full = (socbushandler_wr_lock_counter == 8'd255);
assign socbushandler_wr_lock_empty = (socbushandler_wr_lock_counter == 1'd0);
assign socbushandler_wr_lock_stall = ((cramsoc_aw_valid & cramsoc_aw_ready) & socbushandler_wr_lock_full);
assign socbushandler_rd_lock_full = (socbushandler_rd_lock_counter == 8'd255);
assign socbushandler_rd_lock_empty = (socbushandler_rd_lock_counter == 1'd0);
assign socbushandler_rd_lock_stall = ((cramsoc_ar_valid & cramsoc_ar_ready) & socbushandler_rd_lock_full);
always @(*) begin
    cramsoc_vexriscvaxi_reset_mux <= 32'd1610612736;
    if (cramsoc_trimming_reset_ena) begin
        cramsoc_vexriscvaxi_reset_mux <= cramsoc_trimming_reset;
    end else begin
        cramsoc_vexriscvaxi_reset_mux <= cramsoc_vexriscvaxi;
    end
end
assign cramsoc_zero_trigger = (cramsoc_value == 1'd0);
assign cramsoc_zero0 = cramsoc_zero_status;
assign cramsoc_zero1 = cramsoc_zero_pending;
always @(*) begin
    cramsoc_zero_clear <= 1'd0;
    if ((cramsoc_pending_re & cramsoc_pending_r)) begin
        cramsoc_zero_clear <= 1'd1;
    end
end
assign cramsoc_irq = (cramsoc_pending_status & cramsoc_enable_storage);
assign cramsoc_zero_status = cramsoc_zero_trigger;
assign status = latched_value;
always @(*) begin
    coreuser_coreuser_2bit <= 2'd0;
    if ((cramsoc_satp_asid == {1'd0, coreuser_lut01})) begin
        coreuser_coreuser_2bit <= coreuser_user01;
    end else begin
        if ((cramsoc_satp_asid == {1'd0, coreuser_lut11})) begin
            coreuser_coreuser_2bit <= coreuser_user11;
        end else begin
            if ((cramsoc_satp_asid == {1'd0, coreuser_lut21})) begin
                coreuser_coreuser_2bit <= coreuser_user21;
            end else begin
                if ((cramsoc_satp_asid == {1'd0, coreuser_lut31})) begin
                    coreuser_coreuser_2bit <= coreuser_user31;
                end else begin
                    if ((cramsoc_satp_asid == {1'd0, coreuser_lut41})) begin
                        coreuser_coreuser_2bit <= coreuser_user41;
                    end else begin
                        if ((cramsoc_satp_asid == {1'd0, coreuser_lut51})) begin
                            coreuser_coreuser_2bit <= coreuser_user51;
                        end else begin
                            if ((cramsoc_satp_asid == {1'd0, coreuser_lut61})) begin
                                coreuser_coreuser_2bit <= coreuser_user61;
                            end else begin
                                if ((cramsoc_satp_asid == {1'd0, coreuser_lut71})) begin
                                    coreuser_coreuser_2bit <= coreuser_user71;
                                end else begin
                                    coreuser_coreuser_2bit <= coreuser_user_default;
                                end
                            end
                        end
                    end
                end
            end
        end
    end
end
always @(*) begin
    coreuser_coreuser_4bit <= 4'd0;
    if (coreuser_enable1) begin
        case (coreuser_coreuser_2bit)
            1'd0: begin
                coreuser_coreuser_4bit <= 1'd1;
            end
            1'd1: begin
                coreuser_coreuser_4bit <= 2'd2;
            end
            2'd2: begin
                coreuser_coreuser_4bit <= 3'd4;
            end
            2'd3: begin
                coreuser_coreuser_4bit <= 4'd8;
            end
        endcase
    end else begin
        case (default_user)
            1'd0: begin
                coreuser_coreuser_4bit <= 1'd1;
            end
            1'd1: begin
                coreuser_coreuser_4bit <= 2'd2;
            end
            2'd2: begin
                coreuser_coreuser_4bit <= 3'd4;
            end
            2'd3: begin
                coreuser_coreuser_4bit <= 4'd8;
            end
        endcase
    end
end
assign irqarray0_interrupts = irq_remap0;
assign irqarray0_mdmairq_dupe0 = irqarray0_eventsourceflex0_status;
assign irqarray0_mdmairq_dupe1 = irqarray0_eventsourceflex0_pending;
always @(*) begin
    irqarray0_eventsourceflex0_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[0])) begin
        irqarray0_eventsourceflex0_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s10 = irqarray0_eventsourceflex1_status;
assign irqarray0_nc_b0s11 = irqarray0_eventsourceflex1_pending;
always @(*) begin
    irqarray0_eventsourceflex1_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[1])) begin
        irqarray0_eventsourceflex1_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s20 = irqarray0_eventsourceflex2_status;
assign irqarray0_nc_b0s21 = irqarray0_eventsourceflex2_pending;
always @(*) begin
    irqarray0_eventsourceflex2_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[2])) begin
        irqarray0_eventsourceflex2_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s30 = irqarray0_eventsourceflex3_status;
assign irqarray0_nc_b0s31 = irqarray0_eventsourceflex3_pending;
always @(*) begin
    irqarray0_eventsourceflex3_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[3])) begin
        irqarray0_eventsourceflex3_clear <= 1'd1;
    end
end
assign irqarray0_pioirq0_dupe0 = irqarray0_eventsourceflex4_status;
assign irqarray0_pioirq0_dupe1 = irqarray0_eventsourceflex4_pending;
always @(*) begin
    irqarray0_eventsourceflex4_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[4])) begin
        irqarray0_eventsourceflex4_clear <= 1'd1;
    end
end
assign irqarray0_pioirq1_dupe0 = irqarray0_eventsourceflex5_status;
assign irqarray0_pioirq1_dupe1 = irqarray0_eventsourceflex5_pending;
always @(*) begin
    irqarray0_eventsourceflex5_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[5])) begin
        irqarray0_eventsourceflex5_clear <= 1'd1;
    end
end
assign irqarray0_pioirq2_dupe0 = irqarray0_eventsourceflex6_status;
assign irqarray0_pioirq2_dupe1 = irqarray0_eventsourceflex6_pending;
always @(*) begin
    irqarray0_eventsourceflex6_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[6])) begin
        irqarray0_eventsourceflex6_clear <= 1'd1;
    end
end
assign irqarray0_pioirq3_dupe0 = irqarray0_eventsourceflex7_status;
assign irqarray0_pioirq3_dupe1 = irqarray0_eventsourceflex7_pending;
always @(*) begin
    irqarray0_eventsourceflex7_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[7])) begin
        irqarray0_eventsourceflex7_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s80 = irqarray0_eventsourceflex8_status;
assign irqarray0_nc_b0s81 = irqarray0_eventsourceflex8_pending;
always @(*) begin
    irqarray0_eventsourceflex8_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[8])) begin
        irqarray0_eventsourceflex8_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s90 = irqarray0_eventsourceflex9_status;
assign irqarray0_nc_b0s91 = irqarray0_eventsourceflex9_pending;
always @(*) begin
    irqarray0_eventsourceflex9_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[9])) begin
        irqarray0_eventsourceflex9_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s100 = irqarray0_eventsourceflex10_status;
assign irqarray0_nc_b0s101 = irqarray0_eventsourceflex10_pending;
always @(*) begin
    irqarray0_eventsourceflex10_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[10])) begin
        irqarray0_eventsourceflex10_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s110 = irqarray0_eventsourceflex11_status;
assign irqarray0_nc_b0s111 = irqarray0_eventsourceflex11_pending;
always @(*) begin
    irqarray0_eventsourceflex11_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[11])) begin
        irqarray0_eventsourceflex11_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s120 = irqarray0_eventsourceflex12_status;
assign irqarray0_nc_b0s121 = irqarray0_eventsourceflex12_pending;
always @(*) begin
    irqarray0_eventsourceflex12_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[12])) begin
        irqarray0_eventsourceflex12_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s130 = irqarray0_eventsourceflex13_status;
assign irqarray0_nc_b0s131 = irqarray0_eventsourceflex13_pending;
always @(*) begin
    irqarray0_eventsourceflex13_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[13])) begin
        irqarray0_eventsourceflex13_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s140 = irqarray0_eventsourceflex14_status;
assign irqarray0_nc_b0s141 = irqarray0_eventsourceflex14_pending;
always @(*) begin
    irqarray0_eventsourceflex14_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[14])) begin
        irqarray0_eventsourceflex14_clear <= 1'd1;
    end
end
assign irqarray0_nc_b0s150 = irqarray0_eventsourceflex15_status;
assign irqarray0_nc_b0s151 = irqarray0_eventsourceflex15_pending;
always @(*) begin
    irqarray0_eventsourceflex15_clear <= 1'd0;
    if ((irqarray0_pending_re & irqarray0_pending_r[15])) begin
        irqarray0_eventsourceflex15_clear <= 1'd1;
    end
end
assign irqarray0_irq = ((((((((((((((((irqarray0_pending_status[0] & irqarray0_enable_storage[0]) | (irqarray0_pending_status[1] & irqarray0_enable_storage[1])) | (irqarray0_pending_status[2] & irqarray0_enable_storage[2])) | (irqarray0_pending_status[3] & irqarray0_enable_storage[3])) | (irqarray0_pending_status[4] & irqarray0_enable_storage[4])) | (irqarray0_pending_status[5] & irqarray0_enable_storage[5])) | (irqarray0_pending_status[6] & irqarray0_enable_storage[6])) | (irqarray0_pending_status[7] & irqarray0_enable_storage[7])) | (irqarray0_pending_status[8] & irqarray0_enable_storage[8])) | (irqarray0_pending_status[9] & irqarray0_enable_storage[9])) | (irqarray0_pending_status[10] & irqarray0_enable_storage[10])) | (irqarray0_pending_status[11] & irqarray0_enable_storage[11])) | (irqarray0_pending_status[12] & irqarray0_enable_storage[12])) | (irqarray0_pending_status[13] & irqarray0_enable_storage[13])) | (irqarray0_pending_status[14] & irqarray0_enable_storage[14])) | (irqarray0_pending_status[15] & irqarray0_enable_storage[15]));
always @(*) begin
    irqarray0_eventsourceflex0_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[0]) begin
        if (irqarray0_rising[0]) begin
            irqarray0_eventsourceflex0_trigger_filtered <= (irqarray0_interrupts[0] & (~irqarray0_eventsourceflex0_trigger_d));
        end else begin
            irqarray0_eventsourceflex0_trigger_filtered <= ((~irqarray0_interrupts[0]) & irqarray0_eventsourceflex0_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex0_trigger_filtered <= irqarray0_interrupts[0];
    end
end
assign irqarray0_eventsourceflex0_status = (irqarray0_interrupts[0] | irqarray0_trigger[0]);
always @(*) begin
    irqarray0_eventsourceflex1_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[1]) begin
        if (irqarray0_rising[1]) begin
            irqarray0_eventsourceflex1_trigger_filtered <= (irqarray0_interrupts[1] & (~irqarray0_eventsourceflex1_trigger_d));
        end else begin
            irqarray0_eventsourceflex1_trigger_filtered <= ((~irqarray0_interrupts[1]) & irqarray0_eventsourceflex1_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex1_trigger_filtered <= irqarray0_interrupts[1];
    end
end
assign irqarray0_eventsourceflex1_status = (irqarray0_interrupts[1] | irqarray0_trigger[1]);
always @(*) begin
    irqarray0_eventsourceflex2_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[2]) begin
        if (irqarray0_rising[2]) begin
            irqarray0_eventsourceflex2_trigger_filtered <= (irqarray0_interrupts[2] & (~irqarray0_eventsourceflex2_trigger_d));
        end else begin
            irqarray0_eventsourceflex2_trigger_filtered <= ((~irqarray0_interrupts[2]) & irqarray0_eventsourceflex2_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex2_trigger_filtered <= irqarray0_interrupts[2];
    end
end
assign irqarray0_eventsourceflex2_status = (irqarray0_interrupts[2] | irqarray0_trigger[2]);
always @(*) begin
    irqarray0_eventsourceflex3_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[3]) begin
        if (irqarray0_rising[3]) begin
            irqarray0_eventsourceflex3_trigger_filtered <= (irqarray0_interrupts[3] & (~irqarray0_eventsourceflex3_trigger_d));
        end else begin
            irqarray0_eventsourceflex3_trigger_filtered <= ((~irqarray0_interrupts[3]) & irqarray0_eventsourceflex3_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex3_trigger_filtered <= irqarray0_interrupts[3];
    end
end
assign irqarray0_eventsourceflex3_status = (irqarray0_interrupts[3] | irqarray0_trigger[3]);
always @(*) begin
    irqarray0_eventsourceflex4_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[4]) begin
        if (irqarray0_rising[4]) begin
            irqarray0_eventsourceflex4_trigger_filtered <= (irqarray0_interrupts[4] & (~irqarray0_eventsourceflex4_trigger_d));
        end else begin
            irqarray0_eventsourceflex4_trigger_filtered <= ((~irqarray0_interrupts[4]) & irqarray0_eventsourceflex4_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex4_trigger_filtered <= irqarray0_interrupts[4];
    end
end
assign irqarray0_eventsourceflex4_status = (irqarray0_interrupts[4] | irqarray0_trigger[4]);
always @(*) begin
    irqarray0_eventsourceflex5_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[5]) begin
        if (irqarray0_rising[5]) begin
            irqarray0_eventsourceflex5_trigger_filtered <= (irqarray0_interrupts[5] & (~irqarray0_eventsourceflex5_trigger_d));
        end else begin
            irqarray0_eventsourceflex5_trigger_filtered <= ((~irqarray0_interrupts[5]) & irqarray0_eventsourceflex5_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex5_trigger_filtered <= irqarray0_interrupts[5];
    end
end
assign irqarray0_eventsourceflex5_status = (irqarray0_interrupts[5] | irqarray0_trigger[5]);
always @(*) begin
    irqarray0_eventsourceflex6_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[6]) begin
        if (irqarray0_rising[6]) begin
            irqarray0_eventsourceflex6_trigger_filtered <= (irqarray0_interrupts[6] & (~irqarray0_eventsourceflex6_trigger_d));
        end else begin
            irqarray0_eventsourceflex6_trigger_filtered <= ((~irqarray0_interrupts[6]) & irqarray0_eventsourceflex6_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex6_trigger_filtered <= irqarray0_interrupts[6];
    end
end
assign irqarray0_eventsourceflex6_status = (irqarray0_interrupts[6] | irqarray0_trigger[6]);
always @(*) begin
    irqarray0_eventsourceflex7_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[7]) begin
        if (irqarray0_rising[7]) begin
            irqarray0_eventsourceflex7_trigger_filtered <= (irqarray0_interrupts[7] & (~irqarray0_eventsourceflex7_trigger_d));
        end else begin
            irqarray0_eventsourceflex7_trigger_filtered <= ((~irqarray0_interrupts[7]) & irqarray0_eventsourceflex7_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex7_trigger_filtered <= irqarray0_interrupts[7];
    end
end
assign irqarray0_eventsourceflex7_status = (irqarray0_interrupts[7] | irqarray0_trigger[7]);
always @(*) begin
    irqarray0_eventsourceflex8_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[8]) begin
        if (irqarray0_rising[8]) begin
            irqarray0_eventsourceflex8_trigger_filtered <= (irqarray0_interrupts[8] & (~irqarray0_eventsourceflex8_trigger_d));
        end else begin
            irqarray0_eventsourceflex8_trigger_filtered <= ((~irqarray0_interrupts[8]) & irqarray0_eventsourceflex8_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex8_trigger_filtered <= irqarray0_interrupts[8];
    end
end
assign irqarray0_eventsourceflex8_status = (irqarray0_interrupts[8] | irqarray0_trigger[8]);
always @(*) begin
    irqarray0_eventsourceflex9_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[9]) begin
        if (irqarray0_rising[9]) begin
            irqarray0_eventsourceflex9_trigger_filtered <= (irqarray0_interrupts[9] & (~irqarray0_eventsourceflex9_trigger_d));
        end else begin
            irqarray0_eventsourceflex9_trigger_filtered <= ((~irqarray0_interrupts[9]) & irqarray0_eventsourceflex9_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex9_trigger_filtered <= irqarray0_interrupts[9];
    end
end
assign irqarray0_eventsourceflex9_status = (irqarray0_interrupts[9] | irqarray0_trigger[9]);
always @(*) begin
    irqarray0_eventsourceflex10_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[10]) begin
        if (irqarray0_rising[10]) begin
            irqarray0_eventsourceflex10_trigger_filtered <= (irqarray0_interrupts[10] & (~irqarray0_eventsourceflex10_trigger_d));
        end else begin
            irqarray0_eventsourceflex10_trigger_filtered <= ((~irqarray0_interrupts[10]) & irqarray0_eventsourceflex10_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex10_trigger_filtered <= irqarray0_interrupts[10];
    end
end
assign irqarray0_eventsourceflex10_status = (irqarray0_interrupts[10] | irqarray0_trigger[10]);
always @(*) begin
    irqarray0_eventsourceflex11_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[11]) begin
        if (irqarray0_rising[11]) begin
            irqarray0_eventsourceflex11_trigger_filtered <= (irqarray0_interrupts[11] & (~irqarray0_eventsourceflex11_trigger_d));
        end else begin
            irqarray0_eventsourceflex11_trigger_filtered <= ((~irqarray0_interrupts[11]) & irqarray0_eventsourceflex11_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex11_trigger_filtered <= irqarray0_interrupts[11];
    end
end
assign irqarray0_eventsourceflex11_status = (irqarray0_interrupts[11] | irqarray0_trigger[11]);
always @(*) begin
    irqarray0_eventsourceflex12_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[12]) begin
        if (irqarray0_rising[12]) begin
            irqarray0_eventsourceflex12_trigger_filtered <= (irqarray0_interrupts[12] & (~irqarray0_eventsourceflex12_trigger_d));
        end else begin
            irqarray0_eventsourceflex12_trigger_filtered <= ((~irqarray0_interrupts[12]) & irqarray0_eventsourceflex12_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex12_trigger_filtered <= irqarray0_interrupts[12];
    end
end
assign irqarray0_eventsourceflex12_status = (irqarray0_interrupts[12] | irqarray0_trigger[12]);
always @(*) begin
    irqarray0_eventsourceflex13_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[13]) begin
        if (irqarray0_rising[13]) begin
            irqarray0_eventsourceflex13_trigger_filtered <= (irqarray0_interrupts[13] & (~irqarray0_eventsourceflex13_trigger_d));
        end else begin
            irqarray0_eventsourceflex13_trigger_filtered <= ((~irqarray0_interrupts[13]) & irqarray0_eventsourceflex13_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex13_trigger_filtered <= irqarray0_interrupts[13];
    end
end
assign irqarray0_eventsourceflex13_status = (irqarray0_interrupts[13] | irqarray0_trigger[13]);
always @(*) begin
    irqarray0_eventsourceflex14_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[14]) begin
        if (irqarray0_rising[14]) begin
            irqarray0_eventsourceflex14_trigger_filtered <= (irqarray0_interrupts[14] & (~irqarray0_eventsourceflex14_trigger_d));
        end else begin
            irqarray0_eventsourceflex14_trigger_filtered <= ((~irqarray0_interrupts[14]) & irqarray0_eventsourceflex14_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex14_trigger_filtered <= irqarray0_interrupts[14];
    end
end
assign irqarray0_eventsourceflex14_status = (irqarray0_interrupts[14] | irqarray0_trigger[14]);
always @(*) begin
    irqarray0_eventsourceflex15_trigger_filtered <= 1'd0;
    if (irqarray0_use_edge[15]) begin
        if (irqarray0_rising[15]) begin
            irqarray0_eventsourceflex15_trigger_filtered <= (irqarray0_interrupts[15] & (~irqarray0_eventsourceflex15_trigger_d));
        end else begin
            irqarray0_eventsourceflex15_trigger_filtered <= ((~irqarray0_interrupts[15]) & irqarray0_eventsourceflex15_trigger_d);
        end
    end else begin
        irqarray0_eventsourceflex15_trigger_filtered <= irqarray0_interrupts[15];
    end
end
assign irqarray0_eventsourceflex15_status = (irqarray0_interrupts[15] | irqarray0_trigger[15]);
assign irqarray1_interrupts = irq_remap1;
assign irqarray1_usbc_dupe0 = irqarray1_eventsourceflex16_status;
assign irqarray1_usbc_dupe1 = irqarray1_eventsourceflex16_pending;
always @(*) begin
    irqarray1_eventsourceflex16_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[0])) begin
        irqarray1_eventsourceflex16_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s10 = irqarray1_eventsourceflex17_status;
assign irqarray1_nc_b1s11 = irqarray1_eventsourceflex17_pending;
always @(*) begin
    irqarray1_eventsourceflex17_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[1])) begin
        irqarray1_eventsourceflex17_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s20 = irqarray1_eventsourceflex18_status;
assign irqarray1_nc_b1s21 = irqarray1_eventsourceflex18_pending;
always @(*) begin
    irqarray1_eventsourceflex18_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[2])) begin
        irqarray1_eventsourceflex18_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s30 = irqarray1_eventsourceflex19_status;
assign irqarray1_nc_b1s31 = irqarray1_eventsourceflex19_pending;
always @(*) begin
    irqarray1_eventsourceflex19_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[3])) begin
        irqarray1_eventsourceflex19_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s40 = irqarray1_eventsourceflex20_status;
assign irqarray1_nc_b1s41 = irqarray1_eventsourceflex20_pending;
always @(*) begin
    irqarray1_eventsourceflex20_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[4])) begin
        irqarray1_eventsourceflex20_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s50 = irqarray1_eventsourceflex21_status;
assign irqarray1_nc_b1s51 = irqarray1_eventsourceflex21_pending;
always @(*) begin
    irqarray1_eventsourceflex21_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[5])) begin
        irqarray1_eventsourceflex21_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s60 = irqarray1_eventsourceflex22_status;
assign irqarray1_nc_b1s61 = irqarray1_eventsourceflex22_pending;
always @(*) begin
    irqarray1_eventsourceflex22_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[6])) begin
        irqarray1_eventsourceflex22_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s70 = irqarray1_eventsourceflex23_status;
assign irqarray1_nc_b1s71 = irqarray1_eventsourceflex23_pending;
always @(*) begin
    irqarray1_eventsourceflex23_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[7])) begin
        irqarray1_eventsourceflex23_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s80 = irqarray1_eventsourceflex24_status;
assign irqarray1_nc_b1s81 = irqarray1_eventsourceflex24_pending;
always @(*) begin
    irqarray1_eventsourceflex24_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[8])) begin
        irqarray1_eventsourceflex24_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s90 = irqarray1_eventsourceflex25_status;
assign irqarray1_nc_b1s91 = irqarray1_eventsourceflex25_pending;
always @(*) begin
    irqarray1_eventsourceflex25_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[9])) begin
        irqarray1_eventsourceflex25_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s100 = irqarray1_eventsourceflex26_status;
assign irqarray1_nc_b1s101 = irqarray1_eventsourceflex26_pending;
always @(*) begin
    irqarray1_eventsourceflex26_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[10])) begin
        irqarray1_eventsourceflex26_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s110 = irqarray1_eventsourceflex27_status;
assign irqarray1_nc_b1s111 = irqarray1_eventsourceflex27_pending;
always @(*) begin
    irqarray1_eventsourceflex27_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[11])) begin
        irqarray1_eventsourceflex27_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s120 = irqarray1_eventsourceflex28_status;
assign irqarray1_nc_b1s121 = irqarray1_eventsourceflex28_pending;
always @(*) begin
    irqarray1_eventsourceflex28_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[12])) begin
        irqarray1_eventsourceflex28_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s130 = irqarray1_eventsourceflex29_status;
assign irqarray1_nc_b1s131 = irqarray1_eventsourceflex29_pending;
always @(*) begin
    irqarray1_eventsourceflex29_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[13])) begin
        irqarray1_eventsourceflex29_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s140 = irqarray1_eventsourceflex30_status;
assign irqarray1_nc_b1s141 = irqarray1_eventsourceflex30_pending;
always @(*) begin
    irqarray1_eventsourceflex30_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[14])) begin
        irqarray1_eventsourceflex30_clear <= 1'd1;
    end
end
assign irqarray1_nc_b1s150 = irqarray1_eventsourceflex31_status;
assign irqarray1_nc_b1s151 = irqarray1_eventsourceflex31_pending;
always @(*) begin
    irqarray1_eventsourceflex31_clear <= 1'd0;
    if ((irqarray1_pending_re & irqarray1_pending_r[15])) begin
        irqarray1_eventsourceflex31_clear <= 1'd1;
    end
end
assign irqarray1_irq = ((((((((((((((((irqarray1_pending_status[0] & irqarray1_enable_storage[0]) | (irqarray1_pending_status[1] & irqarray1_enable_storage[1])) | (irqarray1_pending_status[2] & irqarray1_enable_storage[2])) | (irqarray1_pending_status[3] & irqarray1_enable_storage[3])) | (irqarray1_pending_status[4] & irqarray1_enable_storage[4])) | (irqarray1_pending_status[5] & irqarray1_enable_storage[5])) | (irqarray1_pending_status[6] & irqarray1_enable_storage[6])) | (irqarray1_pending_status[7] & irqarray1_enable_storage[7])) | (irqarray1_pending_status[8] & irqarray1_enable_storage[8])) | (irqarray1_pending_status[9] & irqarray1_enable_storage[9])) | (irqarray1_pending_status[10] & irqarray1_enable_storage[10])) | (irqarray1_pending_status[11] & irqarray1_enable_storage[11])) | (irqarray1_pending_status[12] & irqarray1_enable_storage[12])) | (irqarray1_pending_status[13] & irqarray1_enable_storage[13])) | (irqarray1_pending_status[14] & irqarray1_enable_storage[14])) | (irqarray1_pending_status[15] & irqarray1_enable_storage[15]));
always @(*) begin
    irqarray1_eventsourceflex16_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[0]) begin
        if (irqarray1_rising[0]) begin
            irqarray1_eventsourceflex16_trigger_filtered <= (irqarray1_interrupts[0] & (~irqarray1_eventsourceflex16_trigger_d));
        end else begin
            irqarray1_eventsourceflex16_trigger_filtered <= ((~irqarray1_interrupts[0]) & irqarray1_eventsourceflex16_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex16_trigger_filtered <= irqarray1_interrupts[0];
    end
end
assign irqarray1_eventsourceflex16_status = (irqarray1_interrupts[0] | irqarray1_trigger[0]);
always @(*) begin
    irqarray1_eventsourceflex17_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[1]) begin
        if (irqarray1_rising[1]) begin
            irqarray1_eventsourceflex17_trigger_filtered <= (irqarray1_interrupts[1] & (~irqarray1_eventsourceflex17_trigger_d));
        end else begin
            irqarray1_eventsourceflex17_trigger_filtered <= ((~irqarray1_interrupts[1]) & irqarray1_eventsourceflex17_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex17_trigger_filtered <= irqarray1_interrupts[1];
    end
end
assign irqarray1_eventsourceflex17_status = (irqarray1_interrupts[1] | irqarray1_trigger[1]);
always @(*) begin
    irqarray1_eventsourceflex18_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[2]) begin
        if (irqarray1_rising[2]) begin
            irqarray1_eventsourceflex18_trigger_filtered <= (irqarray1_interrupts[2] & (~irqarray1_eventsourceflex18_trigger_d));
        end else begin
            irqarray1_eventsourceflex18_trigger_filtered <= ((~irqarray1_interrupts[2]) & irqarray1_eventsourceflex18_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex18_trigger_filtered <= irqarray1_interrupts[2];
    end
end
assign irqarray1_eventsourceflex18_status = (irqarray1_interrupts[2] | irqarray1_trigger[2]);
always @(*) begin
    irqarray1_eventsourceflex19_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[3]) begin
        if (irqarray1_rising[3]) begin
            irqarray1_eventsourceflex19_trigger_filtered <= (irqarray1_interrupts[3] & (~irqarray1_eventsourceflex19_trigger_d));
        end else begin
            irqarray1_eventsourceflex19_trigger_filtered <= ((~irqarray1_interrupts[3]) & irqarray1_eventsourceflex19_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex19_trigger_filtered <= irqarray1_interrupts[3];
    end
end
assign irqarray1_eventsourceflex19_status = (irqarray1_interrupts[3] | irqarray1_trigger[3]);
always @(*) begin
    irqarray1_eventsourceflex20_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[4]) begin
        if (irqarray1_rising[4]) begin
            irqarray1_eventsourceflex20_trigger_filtered <= (irqarray1_interrupts[4] & (~irqarray1_eventsourceflex20_trigger_d));
        end else begin
            irqarray1_eventsourceflex20_trigger_filtered <= ((~irqarray1_interrupts[4]) & irqarray1_eventsourceflex20_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex20_trigger_filtered <= irqarray1_interrupts[4];
    end
end
assign irqarray1_eventsourceflex20_status = (irqarray1_interrupts[4] | irqarray1_trigger[4]);
always @(*) begin
    irqarray1_eventsourceflex21_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[5]) begin
        if (irqarray1_rising[5]) begin
            irqarray1_eventsourceflex21_trigger_filtered <= (irqarray1_interrupts[5] & (~irqarray1_eventsourceflex21_trigger_d));
        end else begin
            irqarray1_eventsourceflex21_trigger_filtered <= ((~irqarray1_interrupts[5]) & irqarray1_eventsourceflex21_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex21_trigger_filtered <= irqarray1_interrupts[5];
    end
end
assign irqarray1_eventsourceflex21_status = (irqarray1_interrupts[5] | irqarray1_trigger[5]);
always @(*) begin
    irqarray1_eventsourceflex22_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[6]) begin
        if (irqarray1_rising[6]) begin
            irqarray1_eventsourceflex22_trigger_filtered <= (irqarray1_interrupts[6] & (~irqarray1_eventsourceflex22_trigger_d));
        end else begin
            irqarray1_eventsourceflex22_trigger_filtered <= ((~irqarray1_interrupts[6]) & irqarray1_eventsourceflex22_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex22_trigger_filtered <= irqarray1_interrupts[6];
    end
end
assign irqarray1_eventsourceflex22_status = (irqarray1_interrupts[6] | irqarray1_trigger[6]);
always @(*) begin
    irqarray1_eventsourceflex23_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[7]) begin
        if (irqarray1_rising[7]) begin
            irqarray1_eventsourceflex23_trigger_filtered <= (irqarray1_interrupts[7] & (~irqarray1_eventsourceflex23_trigger_d));
        end else begin
            irqarray1_eventsourceflex23_trigger_filtered <= ((~irqarray1_interrupts[7]) & irqarray1_eventsourceflex23_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex23_trigger_filtered <= irqarray1_interrupts[7];
    end
end
assign irqarray1_eventsourceflex23_status = (irqarray1_interrupts[7] | irqarray1_trigger[7]);
always @(*) begin
    irqarray1_eventsourceflex24_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[8]) begin
        if (irqarray1_rising[8]) begin
            irqarray1_eventsourceflex24_trigger_filtered <= (irqarray1_interrupts[8] & (~irqarray1_eventsourceflex24_trigger_d));
        end else begin
            irqarray1_eventsourceflex24_trigger_filtered <= ((~irqarray1_interrupts[8]) & irqarray1_eventsourceflex24_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex24_trigger_filtered <= irqarray1_interrupts[8];
    end
end
assign irqarray1_eventsourceflex24_status = (irqarray1_interrupts[8] | irqarray1_trigger[8]);
always @(*) begin
    irqarray1_eventsourceflex25_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[9]) begin
        if (irqarray1_rising[9]) begin
            irqarray1_eventsourceflex25_trigger_filtered <= (irqarray1_interrupts[9] & (~irqarray1_eventsourceflex25_trigger_d));
        end else begin
            irqarray1_eventsourceflex25_trigger_filtered <= ((~irqarray1_interrupts[9]) & irqarray1_eventsourceflex25_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex25_trigger_filtered <= irqarray1_interrupts[9];
    end
end
assign irqarray1_eventsourceflex25_status = (irqarray1_interrupts[9] | irqarray1_trigger[9]);
always @(*) begin
    irqarray1_eventsourceflex26_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[10]) begin
        if (irqarray1_rising[10]) begin
            irqarray1_eventsourceflex26_trigger_filtered <= (irqarray1_interrupts[10] & (~irqarray1_eventsourceflex26_trigger_d));
        end else begin
            irqarray1_eventsourceflex26_trigger_filtered <= ((~irqarray1_interrupts[10]) & irqarray1_eventsourceflex26_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex26_trigger_filtered <= irqarray1_interrupts[10];
    end
end
assign irqarray1_eventsourceflex26_status = (irqarray1_interrupts[10] | irqarray1_trigger[10]);
always @(*) begin
    irqarray1_eventsourceflex27_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[11]) begin
        if (irqarray1_rising[11]) begin
            irqarray1_eventsourceflex27_trigger_filtered <= (irqarray1_interrupts[11] & (~irqarray1_eventsourceflex27_trigger_d));
        end else begin
            irqarray1_eventsourceflex27_trigger_filtered <= ((~irqarray1_interrupts[11]) & irqarray1_eventsourceflex27_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex27_trigger_filtered <= irqarray1_interrupts[11];
    end
end
assign irqarray1_eventsourceflex27_status = (irqarray1_interrupts[11] | irqarray1_trigger[11]);
always @(*) begin
    irqarray1_eventsourceflex28_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[12]) begin
        if (irqarray1_rising[12]) begin
            irqarray1_eventsourceflex28_trigger_filtered <= (irqarray1_interrupts[12] & (~irqarray1_eventsourceflex28_trigger_d));
        end else begin
            irqarray1_eventsourceflex28_trigger_filtered <= ((~irqarray1_interrupts[12]) & irqarray1_eventsourceflex28_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex28_trigger_filtered <= irqarray1_interrupts[12];
    end
end
assign irqarray1_eventsourceflex28_status = (irqarray1_interrupts[12] | irqarray1_trigger[12]);
always @(*) begin
    irqarray1_eventsourceflex29_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[13]) begin
        if (irqarray1_rising[13]) begin
            irqarray1_eventsourceflex29_trigger_filtered <= (irqarray1_interrupts[13] & (~irqarray1_eventsourceflex29_trigger_d));
        end else begin
            irqarray1_eventsourceflex29_trigger_filtered <= ((~irqarray1_interrupts[13]) & irqarray1_eventsourceflex29_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex29_trigger_filtered <= irqarray1_interrupts[13];
    end
end
assign irqarray1_eventsourceflex29_status = (irqarray1_interrupts[13] | irqarray1_trigger[13]);
always @(*) begin
    irqarray1_eventsourceflex30_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[14]) begin
        if (irqarray1_rising[14]) begin
            irqarray1_eventsourceflex30_trigger_filtered <= (irqarray1_interrupts[14] & (~irqarray1_eventsourceflex30_trigger_d));
        end else begin
            irqarray1_eventsourceflex30_trigger_filtered <= ((~irqarray1_interrupts[14]) & irqarray1_eventsourceflex30_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex30_trigger_filtered <= irqarray1_interrupts[14];
    end
end
assign irqarray1_eventsourceflex30_status = (irqarray1_interrupts[14] | irqarray1_trigger[14]);
always @(*) begin
    irqarray1_eventsourceflex31_trigger_filtered <= 1'd0;
    if (irqarray1_use_edge[15]) begin
        if (irqarray1_rising[15]) begin
            irqarray1_eventsourceflex31_trigger_filtered <= (irqarray1_interrupts[15] & (~irqarray1_eventsourceflex31_trigger_d));
        end else begin
            irqarray1_eventsourceflex31_trigger_filtered <= ((~irqarray1_interrupts[15]) & irqarray1_eventsourceflex31_trigger_d);
        end
    end else begin
        irqarray1_eventsourceflex31_trigger_filtered <= irqarray1_interrupts[15];
    end
end
assign irqarray1_eventsourceflex31_status = (irqarray1_interrupts[15] | irqarray1_trigger[15]);
assign irqarray2_interrupts = irq_remap2;
assign irqarray2_qfcirq0 = irqarray2_eventsourceflex32_status;
assign irqarray2_qfcirq1 = irqarray2_eventsourceflex32_pending;
always @(*) begin
    irqarray2_eventsourceflex32_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[0])) begin
        irqarray2_eventsourceflex32_clear <= 1'd1;
    end
end
assign irqarray2_mdmairq0 = irqarray2_eventsourceflex33_status;
assign irqarray2_mdmairq1 = irqarray2_eventsourceflex33_pending;
always @(*) begin
    irqarray2_eventsourceflex33_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[1])) begin
        irqarray2_eventsourceflex33_clear <= 1'd1;
    end
end
assign irqarray2_mbox_irq_available0 = irqarray2_eventsourceflex34_status;
assign irqarray2_mbox_irq_available1 = irqarray2_eventsourceflex34_pending;
always @(*) begin
    irqarray2_eventsourceflex34_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[2])) begin
        irqarray2_eventsourceflex34_clear <= 1'd1;
    end
end
assign irqarray2_mbox_irq_abort_init0 = irqarray2_eventsourceflex35_status;
assign irqarray2_mbox_irq_abort_init1 = irqarray2_eventsourceflex35_pending;
always @(*) begin
    irqarray2_eventsourceflex35_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[3])) begin
        irqarray2_eventsourceflex35_clear <= 1'd1;
    end
end
assign irqarray2_mbox_irq_done0 = irqarray2_eventsourceflex36_status;
assign irqarray2_mbox_irq_done1 = irqarray2_eventsourceflex36_pending;
always @(*) begin
    irqarray2_eventsourceflex36_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[4])) begin
        irqarray2_eventsourceflex36_clear <= 1'd1;
    end
end
assign irqarray2_mbox_irq_error0 = irqarray2_eventsourceflex37_status;
assign irqarray2_mbox_irq_error1 = irqarray2_eventsourceflex37_pending;
always @(*) begin
    irqarray2_eventsourceflex37_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[5])) begin
        irqarray2_eventsourceflex37_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s60 = irqarray2_eventsourceflex38_status;
assign irqarray2_nc_b2s61 = irqarray2_eventsourceflex38_pending;
always @(*) begin
    irqarray2_eventsourceflex38_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[6])) begin
        irqarray2_eventsourceflex38_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s70 = irqarray2_eventsourceflex39_status;
assign irqarray2_nc_b2s71 = irqarray2_eventsourceflex39_pending;
always @(*) begin
    irqarray2_eventsourceflex39_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[7])) begin
        irqarray2_eventsourceflex39_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s80 = irqarray2_eventsourceflex40_status;
assign irqarray2_nc_b2s81 = irqarray2_eventsourceflex40_pending;
always @(*) begin
    irqarray2_eventsourceflex40_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[8])) begin
        irqarray2_eventsourceflex40_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s90 = irqarray2_eventsourceflex41_status;
assign irqarray2_nc_b2s91 = irqarray2_eventsourceflex41_pending;
always @(*) begin
    irqarray2_eventsourceflex41_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[9])) begin
        irqarray2_eventsourceflex41_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s100 = irqarray2_eventsourceflex42_status;
assign irqarray2_nc_b2s101 = irqarray2_eventsourceflex42_pending;
always @(*) begin
    irqarray2_eventsourceflex42_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[10])) begin
        irqarray2_eventsourceflex42_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s110 = irqarray2_eventsourceflex43_status;
assign irqarray2_nc_b2s111 = irqarray2_eventsourceflex43_pending;
always @(*) begin
    irqarray2_eventsourceflex43_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[11])) begin
        irqarray2_eventsourceflex43_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s120 = irqarray2_eventsourceflex44_status;
assign irqarray2_nc_b2s121 = irqarray2_eventsourceflex44_pending;
always @(*) begin
    irqarray2_eventsourceflex44_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[12])) begin
        irqarray2_eventsourceflex44_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s130 = irqarray2_eventsourceflex45_status;
assign irqarray2_nc_b2s131 = irqarray2_eventsourceflex45_pending;
always @(*) begin
    irqarray2_eventsourceflex45_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[13])) begin
        irqarray2_eventsourceflex45_clear <= 1'd1;
    end
end
assign irqarray2_nc_b2s140 = irqarray2_eventsourceflex46_status;
assign irqarray2_nc_b2s141 = irqarray2_eventsourceflex46_pending;
always @(*) begin
    irqarray2_eventsourceflex46_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[14])) begin
        irqarray2_eventsourceflex46_clear <= 1'd1;
    end
end
assign irqarray2_aowkupint0 = irqarray2_eventsourceflex47_status;
assign irqarray2_aowkupint1 = irqarray2_eventsourceflex47_pending;
always @(*) begin
    irqarray2_eventsourceflex47_clear <= 1'd0;
    if ((irqarray2_pending_re & irqarray2_pending_r[15])) begin
        irqarray2_eventsourceflex47_clear <= 1'd1;
    end
end
assign irqarray2_irq = ((((((((((((((((irqarray2_pending_status[0] & irqarray2_enable_storage[0]) | (irqarray2_pending_status[1] & irqarray2_enable_storage[1])) | (irqarray2_pending_status[2] & irqarray2_enable_storage[2])) | (irqarray2_pending_status[3] & irqarray2_enable_storage[3])) | (irqarray2_pending_status[4] & irqarray2_enable_storage[4])) | (irqarray2_pending_status[5] & irqarray2_enable_storage[5])) | (irqarray2_pending_status[6] & irqarray2_enable_storage[6])) | (irqarray2_pending_status[7] & irqarray2_enable_storage[7])) | (irqarray2_pending_status[8] & irqarray2_enable_storage[8])) | (irqarray2_pending_status[9] & irqarray2_enable_storage[9])) | (irqarray2_pending_status[10] & irqarray2_enable_storage[10])) | (irqarray2_pending_status[11] & irqarray2_enable_storage[11])) | (irqarray2_pending_status[12] & irqarray2_enable_storage[12])) | (irqarray2_pending_status[13] & irqarray2_enable_storage[13])) | (irqarray2_pending_status[14] & irqarray2_enable_storage[14])) | (irqarray2_pending_status[15] & irqarray2_enable_storage[15]));
always @(*) begin
    irqarray2_eventsourceflex32_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[0]) begin
        if (irqarray2_rising[0]) begin
            irqarray2_eventsourceflex32_trigger_filtered <= (irqarray2_interrupts[0] & (~irqarray2_eventsourceflex32_trigger_d));
        end else begin
            irqarray2_eventsourceflex32_trigger_filtered <= ((~irqarray2_interrupts[0]) & irqarray2_eventsourceflex32_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex32_trigger_filtered <= irqarray2_interrupts[0];
    end
end
assign irqarray2_eventsourceflex32_status = (irqarray2_interrupts[0] | irqarray2_trigger[0]);
always @(*) begin
    irqarray2_eventsourceflex33_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[1]) begin
        if (irqarray2_rising[1]) begin
            irqarray2_eventsourceflex33_trigger_filtered <= (irqarray2_interrupts[1] & (~irqarray2_eventsourceflex33_trigger_d));
        end else begin
            irqarray2_eventsourceflex33_trigger_filtered <= ((~irqarray2_interrupts[1]) & irqarray2_eventsourceflex33_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex33_trigger_filtered <= irqarray2_interrupts[1];
    end
end
assign irqarray2_eventsourceflex33_status = (irqarray2_interrupts[1] | irqarray2_trigger[1]);
always @(*) begin
    irqarray2_eventsourceflex34_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[2]) begin
        if (irqarray2_rising[2]) begin
            irqarray2_eventsourceflex34_trigger_filtered <= (irqarray2_interrupts[2] & (~irqarray2_eventsourceflex34_trigger_d));
        end else begin
            irqarray2_eventsourceflex34_trigger_filtered <= ((~irqarray2_interrupts[2]) & irqarray2_eventsourceflex34_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex34_trigger_filtered <= irqarray2_interrupts[2];
    end
end
assign irqarray2_eventsourceflex34_status = (irqarray2_interrupts[2] | irqarray2_trigger[2]);
always @(*) begin
    irqarray2_eventsourceflex35_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[3]) begin
        if (irqarray2_rising[3]) begin
            irqarray2_eventsourceflex35_trigger_filtered <= (irqarray2_interrupts[3] & (~irqarray2_eventsourceflex35_trigger_d));
        end else begin
            irqarray2_eventsourceflex35_trigger_filtered <= ((~irqarray2_interrupts[3]) & irqarray2_eventsourceflex35_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex35_trigger_filtered <= irqarray2_interrupts[3];
    end
end
assign irqarray2_eventsourceflex35_status = (irqarray2_interrupts[3] | irqarray2_trigger[3]);
always @(*) begin
    irqarray2_eventsourceflex36_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[4]) begin
        if (irqarray2_rising[4]) begin
            irqarray2_eventsourceflex36_trigger_filtered <= (irqarray2_interrupts[4] & (~irqarray2_eventsourceflex36_trigger_d));
        end else begin
            irqarray2_eventsourceflex36_trigger_filtered <= ((~irqarray2_interrupts[4]) & irqarray2_eventsourceflex36_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex36_trigger_filtered <= irqarray2_interrupts[4];
    end
end
assign irqarray2_eventsourceflex36_status = (irqarray2_interrupts[4] | irqarray2_trigger[4]);
always @(*) begin
    irqarray2_eventsourceflex37_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[5]) begin
        if (irqarray2_rising[5]) begin
            irqarray2_eventsourceflex37_trigger_filtered <= (irqarray2_interrupts[5] & (~irqarray2_eventsourceflex37_trigger_d));
        end else begin
            irqarray2_eventsourceflex37_trigger_filtered <= ((~irqarray2_interrupts[5]) & irqarray2_eventsourceflex37_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex37_trigger_filtered <= irqarray2_interrupts[5];
    end
end
assign irqarray2_eventsourceflex37_status = (irqarray2_interrupts[5] | irqarray2_trigger[5]);
always @(*) begin
    irqarray2_eventsourceflex38_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[6]) begin
        if (irqarray2_rising[6]) begin
            irqarray2_eventsourceflex38_trigger_filtered <= (irqarray2_interrupts[6] & (~irqarray2_eventsourceflex38_trigger_d));
        end else begin
            irqarray2_eventsourceflex38_trigger_filtered <= ((~irqarray2_interrupts[6]) & irqarray2_eventsourceflex38_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex38_trigger_filtered <= irqarray2_interrupts[6];
    end
end
assign irqarray2_eventsourceflex38_status = (irqarray2_interrupts[6] | irqarray2_trigger[6]);
always @(*) begin
    irqarray2_eventsourceflex39_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[7]) begin
        if (irqarray2_rising[7]) begin
            irqarray2_eventsourceflex39_trigger_filtered <= (irqarray2_interrupts[7] & (~irqarray2_eventsourceflex39_trigger_d));
        end else begin
            irqarray2_eventsourceflex39_trigger_filtered <= ((~irqarray2_interrupts[7]) & irqarray2_eventsourceflex39_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex39_trigger_filtered <= irqarray2_interrupts[7];
    end
end
assign irqarray2_eventsourceflex39_status = (irqarray2_interrupts[7] | irqarray2_trigger[7]);
always @(*) begin
    irqarray2_eventsourceflex40_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[8]) begin
        if (irqarray2_rising[8]) begin
            irqarray2_eventsourceflex40_trigger_filtered <= (irqarray2_interrupts[8] & (~irqarray2_eventsourceflex40_trigger_d));
        end else begin
            irqarray2_eventsourceflex40_trigger_filtered <= ((~irqarray2_interrupts[8]) & irqarray2_eventsourceflex40_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex40_trigger_filtered <= irqarray2_interrupts[8];
    end
end
assign irqarray2_eventsourceflex40_status = (irqarray2_interrupts[8] | irqarray2_trigger[8]);
always @(*) begin
    irqarray2_eventsourceflex41_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[9]) begin
        if (irqarray2_rising[9]) begin
            irqarray2_eventsourceflex41_trigger_filtered <= (irqarray2_interrupts[9] & (~irqarray2_eventsourceflex41_trigger_d));
        end else begin
            irqarray2_eventsourceflex41_trigger_filtered <= ((~irqarray2_interrupts[9]) & irqarray2_eventsourceflex41_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex41_trigger_filtered <= irqarray2_interrupts[9];
    end
end
assign irqarray2_eventsourceflex41_status = (irqarray2_interrupts[9] | irqarray2_trigger[9]);
always @(*) begin
    irqarray2_eventsourceflex42_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[10]) begin
        if (irqarray2_rising[10]) begin
            irqarray2_eventsourceflex42_trigger_filtered <= (irqarray2_interrupts[10] & (~irqarray2_eventsourceflex42_trigger_d));
        end else begin
            irqarray2_eventsourceflex42_trigger_filtered <= ((~irqarray2_interrupts[10]) & irqarray2_eventsourceflex42_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex42_trigger_filtered <= irqarray2_interrupts[10];
    end
end
assign irqarray2_eventsourceflex42_status = (irqarray2_interrupts[10] | irqarray2_trigger[10]);
always @(*) begin
    irqarray2_eventsourceflex43_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[11]) begin
        if (irqarray2_rising[11]) begin
            irqarray2_eventsourceflex43_trigger_filtered <= (irqarray2_interrupts[11] & (~irqarray2_eventsourceflex43_trigger_d));
        end else begin
            irqarray2_eventsourceflex43_trigger_filtered <= ((~irqarray2_interrupts[11]) & irqarray2_eventsourceflex43_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex43_trigger_filtered <= irqarray2_interrupts[11];
    end
end
assign irqarray2_eventsourceflex43_status = (irqarray2_interrupts[11] | irqarray2_trigger[11]);
always @(*) begin
    irqarray2_eventsourceflex44_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[12]) begin
        if (irqarray2_rising[12]) begin
            irqarray2_eventsourceflex44_trigger_filtered <= (irqarray2_interrupts[12] & (~irqarray2_eventsourceflex44_trigger_d));
        end else begin
            irqarray2_eventsourceflex44_trigger_filtered <= ((~irqarray2_interrupts[12]) & irqarray2_eventsourceflex44_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex44_trigger_filtered <= irqarray2_interrupts[12];
    end
end
assign irqarray2_eventsourceflex44_status = (irqarray2_interrupts[12] | irqarray2_trigger[12]);
always @(*) begin
    irqarray2_eventsourceflex45_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[13]) begin
        if (irqarray2_rising[13]) begin
            irqarray2_eventsourceflex45_trigger_filtered <= (irqarray2_interrupts[13] & (~irqarray2_eventsourceflex45_trigger_d));
        end else begin
            irqarray2_eventsourceflex45_trigger_filtered <= ((~irqarray2_interrupts[13]) & irqarray2_eventsourceflex45_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex45_trigger_filtered <= irqarray2_interrupts[13];
    end
end
assign irqarray2_eventsourceflex45_status = (irqarray2_interrupts[13] | irqarray2_trigger[13]);
always @(*) begin
    irqarray2_eventsourceflex46_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[14]) begin
        if (irqarray2_rising[14]) begin
            irqarray2_eventsourceflex46_trigger_filtered <= (irqarray2_interrupts[14] & (~irqarray2_eventsourceflex46_trigger_d));
        end else begin
            irqarray2_eventsourceflex46_trigger_filtered <= ((~irqarray2_interrupts[14]) & irqarray2_eventsourceflex46_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex46_trigger_filtered <= irqarray2_interrupts[14];
    end
end
assign irqarray2_eventsourceflex46_status = (irqarray2_interrupts[14] | irqarray2_trigger[14]);
always @(*) begin
    irqarray2_eventsourceflex47_trigger_filtered <= 1'd0;
    if (irqarray2_use_edge[15]) begin
        if (irqarray2_rising[15]) begin
            irqarray2_eventsourceflex47_trigger_filtered <= (irqarray2_interrupts[15] & (~irqarray2_eventsourceflex47_trigger_d));
        end else begin
            irqarray2_eventsourceflex47_trigger_filtered <= ((~irqarray2_interrupts[15]) & irqarray2_eventsourceflex47_trigger_d);
        end
    end else begin
        irqarray2_eventsourceflex47_trigger_filtered <= irqarray2_interrupts[15];
    end
end
assign irqarray2_eventsourceflex47_status = (irqarray2_interrupts[15] | irqarray2_trigger[15]);
assign irqarray3_interrupts = irq_remap3;
assign irqarray3_trng_done0 = irqarray3_eventsourceflex48_status;
assign irqarray3_trng_done1 = irqarray3_eventsourceflex48_pending;
always @(*) begin
    irqarray3_eventsourceflex48_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[0])) begin
        irqarray3_eventsourceflex48_clear <= 1'd1;
    end
end
assign irqarray3_aes_done0 = irqarray3_eventsourceflex49_status;
assign irqarray3_aes_done1 = irqarray3_eventsourceflex49_pending;
always @(*) begin
    irqarray3_eventsourceflex49_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[1])) begin
        irqarray3_eventsourceflex49_clear <= 1'd1;
    end
end
assign irqarray3_pke_done0 = irqarray3_eventsourceflex50_status;
assign irqarray3_pke_done1 = irqarray3_eventsourceflex50_pending;
always @(*) begin
    irqarray3_eventsourceflex50_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[2])) begin
        irqarray3_eventsourceflex50_clear <= 1'd1;
    end
end
assign irqarray3_hash_done0 = irqarray3_eventsourceflex51_status;
assign irqarray3_hash_done1 = irqarray3_eventsourceflex51_pending;
always @(*) begin
    irqarray3_eventsourceflex51_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[3])) begin
        irqarray3_eventsourceflex51_clear <= 1'd1;
    end
end
assign irqarray3_alu_done0 = irqarray3_eventsourceflex52_status;
assign irqarray3_alu_done1 = irqarray3_eventsourceflex52_pending;
always @(*) begin
    irqarray3_eventsourceflex52_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[4])) begin
        irqarray3_eventsourceflex52_clear <= 1'd1;
    end
end
assign irqarray3_sdma_ichdone0 = irqarray3_eventsourceflex53_status;
assign irqarray3_sdma_ichdone1 = irqarray3_eventsourceflex53_pending;
always @(*) begin
    irqarray3_eventsourceflex53_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[5])) begin
        irqarray3_eventsourceflex53_clear <= 1'd1;
    end
end
assign irqarray3_sdma_schdone0 = irqarray3_eventsourceflex54_status;
assign irqarray3_sdma_schdone1 = irqarray3_eventsourceflex54_pending;
always @(*) begin
    irqarray3_eventsourceflex54_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[6])) begin
        irqarray3_eventsourceflex54_clear <= 1'd1;
    end
end
assign irqarray3_sdma_xchdone0 = irqarray3_eventsourceflex55_status;
assign irqarray3_sdma_xchdone1 = irqarray3_eventsourceflex55_pending;
always @(*) begin
    irqarray3_eventsourceflex55_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[7])) begin
        irqarray3_eventsourceflex55_clear <= 1'd1;
    end
end
assign irqarray3_nc_b3s80 = irqarray3_eventsourceflex56_status;
assign irqarray3_nc_b3s81 = irqarray3_eventsourceflex56_pending;
always @(*) begin
    irqarray3_eventsourceflex56_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[8])) begin
        irqarray3_eventsourceflex56_clear <= 1'd1;
    end
end
assign irqarray3_nc_b3s90 = irqarray3_eventsourceflex57_status;
assign irqarray3_nc_b3s91 = irqarray3_eventsourceflex57_pending;
always @(*) begin
    irqarray3_eventsourceflex57_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[9])) begin
        irqarray3_eventsourceflex57_clear <= 1'd1;
    end
end
assign irqarray3_nc_b3s100 = irqarray3_eventsourceflex58_status;
assign irqarray3_nc_b3s101 = irqarray3_eventsourceflex58_pending;
always @(*) begin
    irqarray3_eventsourceflex58_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[10])) begin
        irqarray3_eventsourceflex58_clear <= 1'd1;
    end
end
assign irqarray3_nc_b3s110 = irqarray3_eventsourceflex59_status;
assign irqarray3_nc_b3s111 = irqarray3_eventsourceflex59_pending;
always @(*) begin
    irqarray3_eventsourceflex59_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[11])) begin
        irqarray3_eventsourceflex59_clear <= 1'd1;
    end
end
assign irqarray3_nc_b3s120 = irqarray3_eventsourceflex60_status;
assign irqarray3_nc_b3s121 = irqarray3_eventsourceflex60_pending;
always @(*) begin
    irqarray3_eventsourceflex60_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[12])) begin
        irqarray3_eventsourceflex60_clear <= 1'd1;
    end
end
assign irqarray3_nc_b3s130 = irqarray3_eventsourceflex61_status;
assign irqarray3_nc_b3s131 = irqarray3_eventsourceflex61_pending;
always @(*) begin
    irqarray3_eventsourceflex61_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[13])) begin
        irqarray3_eventsourceflex61_clear <= 1'd1;
    end
end
assign irqarray3_nc_b3s140 = irqarray3_eventsourceflex62_status;
assign irqarray3_nc_b3s141 = irqarray3_eventsourceflex62_pending;
always @(*) begin
    irqarray3_eventsourceflex62_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[14])) begin
        irqarray3_eventsourceflex62_clear <= 1'd1;
    end
end
assign irqarray3_nc_b3s150 = irqarray3_eventsourceflex63_status;
assign irqarray3_nc_b3s151 = irqarray3_eventsourceflex63_pending;
always @(*) begin
    irqarray3_eventsourceflex63_clear <= 1'd0;
    if ((irqarray3_pending_re & irqarray3_pending_r[15])) begin
        irqarray3_eventsourceflex63_clear <= 1'd1;
    end
end
assign irqarray3_irq = ((((((((((((((((irqarray3_pending_status[0] & irqarray3_enable_storage[0]) | (irqarray3_pending_status[1] & irqarray3_enable_storage[1])) | (irqarray3_pending_status[2] & irqarray3_enable_storage[2])) | (irqarray3_pending_status[3] & irqarray3_enable_storage[3])) | (irqarray3_pending_status[4] & irqarray3_enable_storage[4])) | (irqarray3_pending_status[5] & irqarray3_enable_storage[5])) | (irqarray3_pending_status[6] & irqarray3_enable_storage[6])) | (irqarray3_pending_status[7] & irqarray3_enable_storage[7])) | (irqarray3_pending_status[8] & irqarray3_enable_storage[8])) | (irqarray3_pending_status[9] & irqarray3_enable_storage[9])) | (irqarray3_pending_status[10] & irqarray3_enable_storage[10])) | (irqarray3_pending_status[11] & irqarray3_enable_storage[11])) | (irqarray3_pending_status[12] & irqarray3_enable_storage[12])) | (irqarray3_pending_status[13] & irqarray3_enable_storage[13])) | (irqarray3_pending_status[14] & irqarray3_enable_storage[14])) | (irqarray3_pending_status[15] & irqarray3_enable_storage[15]));
always @(*) begin
    irqarray3_eventsourceflex48_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[0]) begin
        if (irqarray3_rising[0]) begin
            irqarray3_eventsourceflex48_trigger_filtered <= (irqarray3_interrupts[0] & (~irqarray3_eventsourceflex48_trigger_d));
        end else begin
            irqarray3_eventsourceflex48_trigger_filtered <= ((~irqarray3_interrupts[0]) & irqarray3_eventsourceflex48_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex48_trigger_filtered <= irqarray3_interrupts[0];
    end
end
assign irqarray3_eventsourceflex48_status = (irqarray3_interrupts[0] | irqarray3_trigger[0]);
always @(*) begin
    irqarray3_eventsourceflex49_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[1]) begin
        if (irqarray3_rising[1]) begin
            irqarray3_eventsourceflex49_trigger_filtered <= (irqarray3_interrupts[1] & (~irqarray3_eventsourceflex49_trigger_d));
        end else begin
            irqarray3_eventsourceflex49_trigger_filtered <= ((~irqarray3_interrupts[1]) & irqarray3_eventsourceflex49_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex49_trigger_filtered <= irqarray3_interrupts[1];
    end
end
assign irqarray3_eventsourceflex49_status = (irqarray3_interrupts[1] | irqarray3_trigger[1]);
always @(*) begin
    irqarray3_eventsourceflex50_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[2]) begin
        if (irqarray3_rising[2]) begin
            irqarray3_eventsourceflex50_trigger_filtered <= (irqarray3_interrupts[2] & (~irqarray3_eventsourceflex50_trigger_d));
        end else begin
            irqarray3_eventsourceflex50_trigger_filtered <= ((~irqarray3_interrupts[2]) & irqarray3_eventsourceflex50_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex50_trigger_filtered <= irqarray3_interrupts[2];
    end
end
assign irqarray3_eventsourceflex50_status = (irqarray3_interrupts[2] | irqarray3_trigger[2]);
always @(*) begin
    irqarray3_eventsourceflex51_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[3]) begin
        if (irqarray3_rising[3]) begin
            irqarray3_eventsourceflex51_trigger_filtered <= (irqarray3_interrupts[3] & (~irqarray3_eventsourceflex51_trigger_d));
        end else begin
            irqarray3_eventsourceflex51_trigger_filtered <= ((~irqarray3_interrupts[3]) & irqarray3_eventsourceflex51_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex51_trigger_filtered <= irqarray3_interrupts[3];
    end
end
assign irqarray3_eventsourceflex51_status = (irqarray3_interrupts[3] | irqarray3_trigger[3]);
always @(*) begin
    irqarray3_eventsourceflex52_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[4]) begin
        if (irqarray3_rising[4]) begin
            irqarray3_eventsourceflex52_trigger_filtered <= (irqarray3_interrupts[4] & (~irqarray3_eventsourceflex52_trigger_d));
        end else begin
            irqarray3_eventsourceflex52_trigger_filtered <= ((~irqarray3_interrupts[4]) & irqarray3_eventsourceflex52_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex52_trigger_filtered <= irqarray3_interrupts[4];
    end
end
assign irqarray3_eventsourceflex52_status = (irqarray3_interrupts[4] | irqarray3_trigger[4]);
always @(*) begin
    irqarray3_eventsourceflex53_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[5]) begin
        if (irqarray3_rising[5]) begin
            irqarray3_eventsourceflex53_trigger_filtered <= (irqarray3_interrupts[5] & (~irqarray3_eventsourceflex53_trigger_d));
        end else begin
            irqarray3_eventsourceflex53_trigger_filtered <= ((~irqarray3_interrupts[5]) & irqarray3_eventsourceflex53_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex53_trigger_filtered <= irqarray3_interrupts[5];
    end
end
assign irqarray3_eventsourceflex53_status = (irqarray3_interrupts[5] | irqarray3_trigger[5]);
always @(*) begin
    irqarray3_eventsourceflex54_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[6]) begin
        if (irqarray3_rising[6]) begin
            irqarray3_eventsourceflex54_trigger_filtered <= (irqarray3_interrupts[6] & (~irqarray3_eventsourceflex54_trigger_d));
        end else begin
            irqarray3_eventsourceflex54_trigger_filtered <= ((~irqarray3_interrupts[6]) & irqarray3_eventsourceflex54_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex54_trigger_filtered <= irqarray3_interrupts[6];
    end
end
assign irqarray3_eventsourceflex54_status = (irqarray3_interrupts[6] | irqarray3_trigger[6]);
always @(*) begin
    irqarray3_eventsourceflex55_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[7]) begin
        if (irqarray3_rising[7]) begin
            irqarray3_eventsourceflex55_trigger_filtered <= (irqarray3_interrupts[7] & (~irqarray3_eventsourceflex55_trigger_d));
        end else begin
            irqarray3_eventsourceflex55_trigger_filtered <= ((~irqarray3_interrupts[7]) & irqarray3_eventsourceflex55_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex55_trigger_filtered <= irqarray3_interrupts[7];
    end
end
assign irqarray3_eventsourceflex55_status = (irqarray3_interrupts[7] | irqarray3_trigger[7]);
always @(*) begin
    irqarray3_eventsourceflex56_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[8]) begin
        if (irqarray3_rising[8]) begin
            irqarray3_eventsourceflex56_trigger_filtered <= (irqarray3_interrupts[8] & (~irqarray3_eventsourceflex56_trigger_d));
        end else begin
            irqarray3_eventsourceflex56_trigger_filtered <= ((~irqarray3_interrupts[8]) & irqarray3_eventsourceflex56_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex56_trigger_filtered <= irqarray3_interrupts[8];
    end
end
assign irqarray3_eventsourceflex56_status = (irqarray3_interrupts[8] | irqarray3_trigger[8]);
always @(*) begin
    irqarray3_eventsourceflex57_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[9]) begin
        if (irqarray3_rising[9]) begin
            irqarray3_eventsourceflex57_trigger_filtered <= (irqarray3_interrupts[9] & (~irqarray3_eventsourceflex57_trigger_d));
        end else begin
            irqarray3_eventsourceflex57_trigger_filtered <= ((~irqarray3_interrupts[9]) & irqarray3_eventsourceflex57_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex57_trigger_filtered <= irqarray3_interrupts[9];
    end
end
assign irqarray3_eventsourceflex57_status = (irqarray3_interrupts[9] | irqarray3_trigger[9]);
always @(*) begin
    irqarray3_eventsourceflex58_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[10]) begin
        if (irqarray3_rising[10]) begin
            irqarray3_eventsourceflex58_trigger_filtered <= (irqarray3_interrupts[10] & (~irqarray3_eventsourceflex58_trigger_d));
        end else begin
            irqarray3_eventsourceflex58_trigger_filtered <= ((~irqarray3_interrupts[10]) & irqarray3_eventsourceflex58_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex58_trigger_filtered <= irqarray3_interrupts[10];
    end
end
assign irqarray3_eventsourceflex58_status = (irqarray3_interrupts[10] | irqarray3_trigger[10]);
always @(*) begin
    irqarray3_eventsourceflex59_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[11]) begin
        if (irqarray3_rising[11]) begin
            irqarray3_eventsourceflex59_trigger_filtered <= (irqarray3_interrupts[11] & (~irqarray3_eventsourceflex59_trigger_d));
        end else begin
            irqarray3_eventsourceflex59_trigger_filtered <= ((~irqarray3_interrupts[11]) & irqarray3_eventsourceflex59_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex59_trigger_filtered <= irqarray3_interrupts[11];
    end
end
assign irqarray3_eventsourceflex59_status = (irqarray3_interrupts[11] | irqarray3_trigger[11]);
always @(*) begin
    irqarray3_eventsourceflex60_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[12]) begin
        if (irqarray3_rising[12]) begin
            irqarray3_eventsourceflex60_trigger_filtered <= (irqarray3_interrupts[12] & (~irqarray3_eventsourceflex60_trigger_d));
        end else begin
            irqarray3_eventsourceflex60_trigger_filtered <= ((~irqarray3_interrupts[12]) & irqarray3_eventsourceflex60_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex60_trigger_filtered <= irqarray3_interrupts[12];
    end
end
assign irqarray3_eventsourceflex60_status = (irqarray3_interrupts[12] | irqarray3_trigger[12]);
always @(*) begin
    irqarray3_eventsourceflex61_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[13]) begin
        if (irqarray3_rising[13]) begin
            irqarray3_eventsourceflex61_trigger_filtered <= (irqarray3_interrupts[13] & (~irqarray3_eventsourceflex61_trigger_d));
        end else begin
            irqarray3_eventsourceflex61_trigger_filtered <= ((~irqarray3_interrupts[13]) & irqarray3_eventsourceflex61_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex61_trigger_filtered <= irqarray3_interrupts[13];
    end
end
assign irqarray3_eventsourceflex61_status = (irqarray3_interrupts[13] | irqarray3_trigger[13]);
always @(*) begin
    irqarray3_eventsourceflex62_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[14]) begin
        if (irqarray3_rising[14]) begin
            irqarray3_eventsourceflex62_trigger_filtered <= (irqarray3_interrupts[14] & (~irqarray3_eventsourceflex62_trigger_d));
        end else begin
            irqarray3_eventsourceflex62_trigger_filtered <= ((~irqarray3_interrupts[14]) & irqarray3_eventsourceflex62_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex62_trigger_filtered <= irqarray3_interrupts[14];
    end
end
assign irqarray3_eventsourceflex62_status = (irqarray3_interrupts[14] | irqarray3_trigger[14]);
always @(*) begin
    irqarray3_eventsourceflex63_trigger_filtered <= 1'd0;
    if (irqarray3_use_edge[15]) begin
        if (irqarray3_rising[15]) begin
            irqarray3_eventsourceflex63_trigger_filtered <= (irqarray3_interrupts[15] & (~irqarray3_eventsourceflex63_trigger_d));
        end else begin
            irqarray3_eventsourceflex63_trigger_filtered <= ((~irqarray3_interrupts[15]) & irqarray3_eventsourceflex63_trigger_d);
        end
    end else begin
        irqarray3_eventsourceflex63_trigger_filtered <= irqarray3_interrupts[15];
    end
end
assign irqarray3_eventsourceflex63_status = (irqarray3_interrupts[15] | irqarray3_trigger[15]);
assign irqarray4_interrupts = irq_remap4;
assign irqarray4_trng_done_dupe0 = irqarray4_eventsourceflex64_status;
assign irqarray4_trng_done_dupe1 = irqarray4_eventsourceflex64_pending;
always @(*) begin
    irqarray4_eventsourceflex64_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[0])) begin
        irqarray4_eventsourceflex64_clear <= 1'd1;
    end
end
assign irqarray4_aes_done_dupe0 = irqarray4_eventsourceflex65_status;
assign irqarray4_aes_done_dupe1 = irqarray4_eventsourceflex65_pending;
always @(*) begin
    irqarray4_eventsourceflex65_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[1])) begin
        irqarray4_eventsourceflex65_clear <= 1'd1;
    end
end
assign irqarray4_pke_done_dupe0 = irqarray4_eventsourceflex66_status;
assign irqarray4_pke_done_dupe1 = irqarray4_eventsourceflex66_pending;
always @(*) begin
    irqarray4_eventsourceflex66_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[2])) begin
        irqarray4_eventsourceflex66_clear <= 1'd1;
    end
end
assign irqarray4_hash_done_dupe0 = irqarray4_eventsourceflex67_status;
assign irqarray4_hash_done_dupe1 = irqarray4_eventsourceflex67_pending;
always @(*) begin
    irqarray4_eventsourceflex67_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[3])) begin
        irqarray4_eventsourceflex67_clear <= 1'd1;
    end
end
assign irqarray4_alu_done_dupe0 = irqarray4_eventsourceflex68_status;
assign irqarray4_alu_done_dupe1 = irqarray4_eventsourceflex68_pending;
always @(*) begin
    irqarray4_eventsourceflex68_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[4])) begin
        irqarray4_eventsourceflex68_clear <= 1'd1;
    end
end
assign irqarray4_sdma_ichdone_dupe0 = irqarray4_eventsourceflex69_status;
assign irqarray4_sdma_ichdone_dupe1 = irqarray4_eventsourceflex69_pending;
always @(*) begin
    irqarray4_eventsourceflex69_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[5])) begin
        irqarray4_eventsourceflex69_clear <= 1'd1;
    end
end
assign irqarray4_sdma_schdone_dupe0 = irqarray4_eventsourceflex70_status;
assign irqarray4_sdma_schdone_dupe1 = irqarray4_eventsourceflex70_pending;
always @(*) begin
    irqarray4_eventsourceflex70_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[6])) begin
        irqarray4_eventsourceflex70_clear <= 1'd1;
    end
end
assign irqarray4_sdma_xchdone_dupe0 = irqarray4_eventsourceflex71_status;
assign irqarray4_sdma_xchdone_dupe1 = irqarray4_eventsourceflex71_pending;
always @(*) begin
    irqarray4_eventsourceflex71_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[7])) begin
        irqarray4_eventsourceflex71_clear <= 1'd1;
    end
end
assign irqarray4_nc_b4s80 = irqarray4_eventsourceflex72_status;
assign irqarray4_nc_b4s81 = irqarray4_eventsourceflex72_pending;
always @(*) begin
    irqarray4_eventsourceflex72_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[8])) begin
        irqarray4_eventsourceflex72_clear <= 1'd1;
    end
end
assign irqarray4_nc_b4s90 = irqarray4_eventsourceflex73_status;
assign irqarray4_nc_b4s91 = irqarray4_eventsourceflex73_pending;
always @(*) begin
    irqarray4_eventsourceflex73_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[9])) begin
        irqarray4_eventsourceflex73_clear <= 1'd1;
    end
end
assign irqarray4_nc_b4s100 = irqarray4_eventsourceflex74_status;
assign irqarray4_nc_b4s101 = irqarray4_eventsourceflex74_pending;
always @(*) begin
    irqarray4_eventsourceflex74_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[10])) begin
        irqarray4_eventsourceflex74_clear <= 1'd1;
    end
end
assign irqarray4_nc_b4s110 = irqarray4_eventsourceflex75_status;
assign irqarray4_nc_b4s111 = irqarray4_eventsourceflex75_pending;
always @(*) begin
    irqarray4_eventsourceflex75_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[11])) begin
        irqarray4_eventsourceflex75_clear <= 1'd1;
    end
end
assign irqarray4_nc_b4s120 = irqarray4_eventsourceflex76_status;
assign irqarray4_nc_b4s121 = irqarray4_eventsourceflex76_pending;
always @(*) begin
    irqarray4_eventsourceflex76_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[12])) begin
        irqarray4_eventsourceflex76_clear <= 1'd1;
    end
end
assign irqarray4_nc_b4s130 = irqarray4_eventsourceflex77_status;
assign irqarray4_nc_b4s131 = irqarray4_eventsourceflex77_pending;
always @(*) begin
    irqarray4_eventsourceflex77_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[13])) begin
        irqarray4_eventsourceflex77_clear <= 1'd1;
    end
end
assign irqarray4_nc_b4s140 = irqarray4_eventsourceflex78_status;
assign irqarray4_nc_b4s141 = irqarray4_eventsourceflex78_pending;
always @(*) begin
    irqarray4_eventsourceflex78_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[14])) begin
        irqarray4_eventsourceflex78_clear <= 1'd1;
    end
end
assign irqarray4_nc_b4s150 = irqarray4_eventsourceflex79_status;
assign irqarray4_nc_b4s151 = irqarray4_eventsourceflex79_pending;
always @(*) begin
    irqarray4_eventsourceflex79_clear <= 1'd0;
    if ((irqarray4_pending_re & irqarray4_pending_r[15])) begin
        irqarray4_eventsourceflex79_clear <= 1'd1;
    end
end
assign irqarray4_irq = ((((((((((((((((irqarray4_pending_status[0] & irqarray4_enable_storage[0]) | (irqarray4_pending_status[1] & irqarray4_enable_storage[1])) | (irqarray4_pending_status[2] & irqarray4_enable_storage[2])) | (irqarray4_pending_status[3] & irqarray4_enable_storage[3])) | (irqarray4_pending_status[4] & irqarray4_enable_storage[4])) | (irqarray4_pending_status[5] & irqarray4_enable_storage[5])) | (irqarray4_pending_status[6] & irqarray4_enable_storage[6])) | (irqarray4_pending_status[7] & irqarray4_enable_storage[7])) | (irqarray4_pending_status[8] & irqarray4_enable_storage[8])) | (irqarray4_pending_status[9] & irqarray4_enable_storage[9])) | (irqarray4_pending_status[10] & irqarray4_enable_storage[10])) | (irqarray4_pending_status[11] & irqarray4_enable_storage[11])) | (irqarray4_pending_status[12] & irqarray4_enable_storage[12])) | (irqarray4_pending_status[13] & irqarray4_enable_storage[13])) | (irqarray4_pending_status[14] & irqarray4_enable_storage[14])) | (irqarray4_pending_status[15] & irqarray4_enable_storage[15]));
always @(*) begin
    irqarray4_eventsourceflex64_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[0]) begin
        if (irqarray4_rising[0]) begin
            irqarray4_eventsourceflex64_trigger_filtered <= (irqarray4_interrupts[0] & (~irqarray4_eventsourceflex64_trigger_d));
        end else begin
            irqarray4_eventsourceflex64_trigger_filtered <= ((~irqarray4_interrupts[0]) & irqarray4_eventsourceflex64_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex64_trigger_filtered <= irqarray4_interrupts[0];
    end
end
assign irqarray4_eventsourceflex64_status = (irqarray4_interrupts[0] | irqarray4_trigger[0]);
always @(*) begin
    irqarray4_eventsourceflex65_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[1]) begin
        if (irqarray4_rising[1]) begin
            irqarray4_eventsourceflex65_trigger_filtered <= (irqarray4_interrupts[1] & (~irqarray4_eventsourceflex65_trigger_d));
        end else begin
            irqarray4_eventsourceflex65_trigger_filtered <= ((~irqarray4_interrupts[1]) & irqarray4_eventsourceflex65_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex65_trigger_filtered <= irqarray4_interrupts[1];
    end
end
assign irqarray4_eventsourceflex65_status = (irqarray4_interrupts[1] | irqarray4_trigger[1]);
always @(*) begin
    irqarray4_eventsourceflex66_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[2]) begin
        if (irqarray4_rising[2]) begin
            irqarray4_eventsourceflex66_trigger_filtered <= (irqarray4_interrupts[2] & (~irqarray4_eventsourceflex66_trigger_d));
        end else begin
            irqarray4_eventsourceflex66_trigger_filtered <= ((~irqarray4_interrupts[2]) & irqarray4_eventsourceflex66_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex66_trigger_filtered <= irqarray4_interrupts[2];
    end
end
assign irqarray4_eventsourceflex66_status = (irqarray4_interrupts[2] | irqarray4_trigger[2]);
always @(*) begin
    irqarray4_eventsourceflex67_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[3]) begin
        if (irqarray4_rising[3]) begin
            irqarray4_eventsourceflex67_trigger_filtered <= (irqarray4_interrupts[3] & (~irqarray4_eventsourceflex67_trigger_d));
        end else begin
            irqarray4_eventsourceflex67_trigger_filtered <= ((~irqarray4_interrupts[3]) & irqarray4_eventsourceflex67_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex67_trigger_filtered <= irqarray4_interrupts[3];
    end
end
assign irqarray4_eventsourceflex67_status = (irqarray4_interrupts[3] | irqarray4_trigger[3]);
always @(*) begin
    irqarray4_eventsourceflex68_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[4]) begin
        if (irqarray4_rising[4]) begin
            irqarray4_eventsourceflex68_trigger_filtered <= (irqarray4_interrupts[4] & (~irqarray4_eventsourceflex68_trigger_d));
        end else begin
            irqarray4_eventsourceflex68_trigger_filtered <= ((~irqarray4_interrupts[4]) & irqarray4_eventsourceflex68_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex68_trigger_filtered <= irqarray4_interrupts[4];
    end
end
assign irqarray4_eventsourceflex68_status = (irqarray4_interrupts[4] | irqarray4_trigger[4]);
always @(*) begin
    irqarray4_eventsourceflex69_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[5]) begin
        if (irqarray4_rising[5]) begin
            irqarray4_eventsourceflex69_trigger_filtered <= (irqarray4_interrupts[5] & (~irqarray4_eventsourceflex69_trigger_d));
        end else begin
            irqarray4_eventsourceflex69_trigger_filtered <= ((~irqarray4_interrupts[5]) & irqarray4_eventsourceflex69_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex69_trigger_filtered <= irqarray4_interrupts[5];
    end
end
assign irqarray4_eventsourceflex69_status = (irqarray4_interrupts[5] | irqarray4_trigger[5]);
always @(*) begin
    irqarray4_eventsourceflex70_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[6]) begin
        if (irqarray4_rising[6]) begin
            irqarray4_eventsourceflex70_trigger_filtered <= (irqarray4_interrupts[6] & (~irqarray4_eventsourceflex70_trigger_d));
        end else begin
            irqarray4_eventsourceflex70_trigger_filtered <= ((~irqarray4_interrupts[6]) & irqarray4_eventsourceflex70_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex70_trigger_filtered <= irqarray4_interrupts[6];
    end
end
assign irqarray4_eventsourceflex70_status = (irqarray4_interrupts[6] | irqarray4_trigger[6]);
always @(*) begin
    irqarray4_eventsourceflex71_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[7]) begin
        if (irqarray4_rising[7]) begin
            irqarray4_eventsourceflex71_trigger_filtered <= (irqarray4_interrupts[7] & (~irqarray4_eventsourceflex71_trigger_d));
        end else begin
            irqarray4_eventsourceflex71_trigger_filtered <= ((~irqarray4_interrupts[7]) & irqarray4_eventsourceflex71_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex71_trigger_filtered <= irqarray4_interrupts[7];
    end
end
assign irqarray4_eventsourceflex71_status = (irqarray4_interrupts[7] | irqarray4_trigger[7]);
always @(*) begin
    irqarray4_eventsourceflex72_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[8]) begin
        if (irqarray4_rising[8]) begin
            irqarray4_eventsourceflex72_trigger_filtered <= (irqarray4_interrupts[8] & (~irqarray4_eventsourceflex72_trigger_d));
        end else begin
            irqarray4_eventsourceflex72_trigger_filtered <= ((~irqarray4_interrupts[8]) & irqarray4_eventsourceflex72_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex72_trigger_filtered <= irqarray4_interrupts[8];
    end
end
assign irqarray4_eventsourceflex72_status = (irqarray4_interrupts[8] | irqarray4_trigger[8]);
always @(*) begin
    irqarray4_eventsourceflex73_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[9]) begin
        if (irqarray4_rising[9]) begin
            irqarray4_eventsourceflex73_trigger_filtered <= (irqarray4_interrupts[9] & (~irqarray4_eventsourceflex73_trigger_d));
        end else begin
            irqarray4_eventsourceflex73_trigger_filtered <= ((~irqarray4_interrupts[9]) & irqarray4_eventsourceflex73_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex73_trigger_filtered <= irqarray4_interrupts[9];
    end
end
assign irqarray4_eventsourceflex73_status = (irqarray4_interrupts[9] | irqarray4_trigger[9]);
always @(*) begin
    irqarray4_eventsourceflex74_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[10]) begin
        if (irqarray4_rising[10]) begin
            irqarray4_eventsourceflex74_trigger_filtered <= (irqarray4_interrupts[10] & (~irqarray4_eventsourceflex74_trigger_d));
        end else begin
            irqarray4_eventsourceflex74_trigger_filtered <= ((~irqarray4_interrupts[10]) & irqarray4_eventsourceflex74_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex74_trigger_filtered <= irqarray4_interrupts[10];
    end
end
assign irqarray4_eventsourceflex74_status = (irqarray4_interrupts[10] | irqarray4_trigger[10]);
always @(*) begin
    irqarray4_eventsourceflex75_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[11]) begin
        if (irqarray4_rising[11]) begin
            irqarray4_eventsourceflex75_trigger_filtered <= (irqarray4_interrupts[11] & (~irqarray4_eventsourceflex75_trigger_d));
        end else begin
            irqarray4_eventsourceflex75_trigger_filtered <= ((~irqarray4_interrupts[11]) & irqarray4_eventsourceflex75_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex75_trigger_filtered <= irqarray4_interrupts[11];
    end
end
assign irqarray4_eventsourceflex75_status = (irqarray4_interrupts[11] | irqarray4_trigger[11]);
always @(*) begin
    irqarray4_eventsourceflex76_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[12]) begin
        if (irqarray4_rising[12]) begin
            irqarray4_eventsourceflex76_trigger_filtered <= (irqarray4_interrupts[12] & (~irqarray4_eventsourceflex76_trigger_d));
        end else begin
            irqarray4_eventsourceflex76_trigger_filtered <= ((~irqarray4_interrupts[12]) & irqarray4_eventsourceflex76_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex76_trigger_filtered <= irqarray4_interrupts[12];
    end
end
assign irqarray4_eventsourceflex76_status = (irqarray4_interrupts[12] | irqarray4_trigger[12]);
always @(*) begin
    irqarray4_eventsourceflex77_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[13]) begin
        if (irqarray4_rising[13]) begin
            irqarray4_eventsourceflex77_trigger_filtered <= (irqarray4_interrupts[13] & (~irqarray4_eventsourceflex77_trigger_d));
        end else begin
            irqarray4_eventsourceflex77_trigger_filtered <= ((~irqarray4_interrupts[13]) & irqarray4_eventsourceflex77_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex77_trigger_filtered <= irqarray4_interrupts[13];
    end
end
assign irqarray4_eventsourceflex77_status = (irqarray4_interrupts[13] | irqarray4_trigger[13]);
always @(*) begin
    irqarray4_eventsourceflex78_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[14]) begin
        if (irqarray4_rising[14]) begin
            irqarray4_eventsourceflex78_trigger_filtered <= (irqarray4_interrupts[14] & (~irqarray4_eventsourceflex78_trigger_d));
        end else begin
            irqarray4_eventsourceflex78_trigger_filtered <= ((~irqarray4_interrupts[14]) & irqarray4_eventsourceflex78_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex78_trigger_filtered <= irqarray4_interrupts[14];
    end
end
assign irqarray4_eventsourceflex78_status = (irqarray4_interrupts[14] | irqarray4_trigger[14]);
always @(*) begin
    irqarray4_eventsourceflex79_trigger_filtered <= 1'd0;
    if (irqarray4_use_edge[15]) begin
        if (irqarray4_rising[15]) begin
            irqarray4_eventsourceflex79_trigger_filtered <= (irqarray4_interrupts[15] & (~irqarray4_eventsourceflex79_trigger_d));
        end else begin
            irqarray4_eventsourceflex79_trigger_filtered <= ((~irqarray4_interrupts[15]) & irqarray4_eventsourceflex79_trigger_d);
        end
    end else begin
        irqarray4_eventsourceflex79_trigger_filtered <= irqarray4_interrupts[15];
    end
end
assign irqarray4_eventsourceflex79_status = (irqarray4_interrupts[15] | irqarray4_trigger[15]);
assign irqarray5_interrupts = irq_remap5;
assign irqarray5_uart0_rx0 = irqarray5_eventsourceflex80_status;
assign irqarray5_uart0_rx1 = irqarray5_eventsourceflex80_pending;
always @(*) begin
    irqarray5_eventsourceflex80_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[0])) begin
        irqarray5_eventsourceflex80_clear <= 1'd1;
    end
end
assign irqarray5_uart0_tx0 = irqarray5_eventsourceflex81_status;
assign irqarray5_uart0_tx1 = irqarray5_eventsourceflex81_pending;
always @(*) begin
    irqarray5_eventsourceflex81_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[1])) begin
        irqarray5_eventsourceflex81_clear <= 1'd1;
    end
end
assign irqarray5_uart0_rx_char0 = irqarray5_eventsourceflex82_status;
assign irqarray5_uart0_rx_char1 = irqarray5_eventsourceflex82_pending;
always @(*) begin
    irqarray5_eventsourceflex82_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[2])) begin
        irqarray5_eventsourceflex82_clear <= 1'd1;
    end
end
assign irqarray5_uart0_err0 = irqarray5_eventsourceflex83_status;
assign irqarray5_uart0_err1 = irqarray5_eventsourceflex83_pending;
always @(*) begin
    irqarray5_eventsourceflex83_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[3])) begin
        irqarray5_eventsourceflex83_clear <= 1'd1;
    end
end
assign irqarray5_uart1_rx0 = irqarray5_eventsourceflex84_status;
assign irqarray5_uart1_rx1 = irqarray5_eventsourceflex84_pending;
always @(*) begin
    irqarray5_eventsourceflex84_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[4])) begin
        irqarray5_eventsourceflex84_clear <= 1'd1;
    end
end
assign irqarray5_uart1_tx0 = irqarray5_eventsourceflex85_status;
assign irqarray5_uart1_tx1 = irqarray5_eventsourceflex85_pending;
always @(*) begin
    irqarray5_eventsourceflex85_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[5])) begin
        irqarray5_eventsourceflex85_clear <= 1'd1;
    end
end
assign irqarray5_uart1_rx_char0 = irqarray5_eventsourceflex86_status;
assign irqarray5_uart1_rx_char1 = irqarray5_eventsourceflex86_pending;
always @(*) begin
    irqarray5_eventsourceflex86_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[6])) begin
        irqarray5_eventsourceflex86_clear <= 1'd1;
    end
end
assign irqarray5_uart1_err0 = irqarray5_eventsourceflex87_status;
assign irqarray5_uart1_err1 = irqarray5_eventsourceflex87_pending;
always @(*) begin
    irqarray5_eventsourceflex87_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[7])) begin
        irqarray5_eventsourceflex87_clear <= 1'd1;
    end
end
assign irqarray5_uart2_rx0 = irqarray5_eventsourceflex88_status;
assign irqarray5_uart2_rx1 = irqarray5_eventsourceflex88_pending;
always @(*) begin
    irqarray5_eventsourceflex88_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[8])) begin
        irqarray5_eventsourceflex88_clear <= 1'd1;
    end
end
assign irqarray5_uart2_tx0 = irqarray5_eventsourceflex89_status;
assign irqarray5_uart2_tx1 = irqarray5_eventsourceflex89_pending;
always @(*) begin
    irqarray5_eventsourceflex89_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[9])) begin
        irqarray5_eventsourceflex89_clear <= 1'd1;
    end
end
assign irqarray5_uart2_rx_char0 = irqarray5_eventsourceflex90_status;
assign irqarray5_uart2_rx_char1 = irqarray5_eventsourceflex90_pending;
always @(*) begin
    irqarray5_eventsourceflex90_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[10])) begin
        irqarray5_eventsourceflex90_clear <= 1'd1;
    end
end
assign irqarray5_uart2_err0 = irqarray5_eventsourceflex91_status;
assign irqarray5_uart2_err1 = irqarray5_eventsourceflex91_pending;
always @(*) begin
    irqarray5_eventsourceflex91_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[11])) begin
        irqarray5_eventsourceflex91_clear <= 1'd1;
    end
end
assign irqarray5_uart3_rx0 = irqarray5_eventsourceflex92_status;
assign irqarray5_uart3_rx1 = irqarray5_eventsourceflex92_pending;
always @(*) begin
    irqarray5_eventsourceflex92_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[12])) begin
        irqarray5_eventsourceflex92_clear <= 1'd1;
    end
end
assign irqarray5_uart3_tx0 = irqarray5_eventsourceflex93_status;
assign irqarray5_uart3_tx1 = irqarray5_eventsourceflex93_pending;
always @(*) begin
    irqarray5_eventsourceflex93_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[13])) begin
        irqarray5_eventsourceflex93_clear <= 1'd1;
    end
end
assign irqarray5_uart3_rx_char0 = irqarray5_eventsourceflex94_status;
assign irqarray5_uart3_rx_char1 = irqarray5_eventsourceflex94_pending;
always @(*) begin
    irqarray5_eventsourceflex94_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[14])) begin
        irqarray5_eventsourceflex94_clear <= 1'd1;
    end
end
assign irqarray5_uart3_err0 = irqarray5_eventsourceflex95_status;
assign irqarray5_uart3_err1 = irqarray5_eventsourceflex95_pending;
always @(*) begin
    irqarray5_eventsourceflex95_clear <= 1'd0;
    if ((irqarray5_pending_re & irqarray5_pending_r[15])) begin
        irqarray5_eventsourceflex95_clear <= 1'd1;
    end
end
assign irqarray5_irq = ((((((((((((((((irqarray5_pending_status[0] & irqarray5_enable_storage[0]) | (irqarray5_pending_status[1] & irqarray5_enable_storage[1])) | (irqarray5_pending_status[2] & irqarray5_enable_storage[2])) | (irqarray5_pending_status[3] & irqarray5_enable_storage[3])) | (irqarray5_pending_status[4] & irqarray5_enable_storage[4])) | (irqarray5_pending_status[5] & irqarray5_enable_storage[5])) | (irqarray5_pending_status[6] & irqarray5_enable_storage[6])) | (irqarray5_pending_status[7] & irqarray5_enable_storage[7])) | (irqarray5_pending_status[8] & irqarray5_enable_storage[8])) | (irqarray5_pending_status[9] & irqarray5_enable_storage[9])) | (irqarray5_pending_status[10] & irqarray5_enable_storage[10])) | (irqarray5_pending_status[11] & irqarray5_enable_storage[11])) | (irqarray5_pending_status[12] & irqarray5_enable_storage[12])) | (irqarray5_pending_status[13] & irqarray5_enable_storage[13])) | (irqarray5_pending_status[14] & irqarray5_enable_storage[14])) | (irqarray5_pending_status[15] & irqarray5_enable_storage[15]));
always @(*) begin
    irqarray5_eventsourceflex80_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[0]) begin
        if (irqarray5_rising[0]) begin
            irqarray5_eventsourceflex80_trigger_filtered <= (irqarray5_interrupts[0] & (~irqarray5_eventsourceflex80_trigger_d));
        end else begin
            irqarray5_eventsourceflex80_trigger_filtered <= ((~irqarray5_interrupts[0]) & irqarray5_eventsourceflex80_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex80_trigger_filtered <= irqarray5_interrupts[0];
    end
end
assign irqarray5_eventsourceflex80_status = (irqarray5_interrupts[0] | irqarray5_trigger[0]);
always @(*) begin
    irqarray5_eventsourceflex81_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[1]) begin
        if (irqarray5_rising[1]) begin
            irqarray5_eventsourceflex81_trigger_filtered <= (irqarray5_interrupts[1] & (~irqarray5_eventsourceflex81_trigger_d));
        end else begin
            irqarray5_eventsourceflex81_trigger_filtered <= ((~irqarray5_interrupts[1]) & irqarray5_eventsourceflex81_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex81_trigger_filtered <= irqarray5_interrupts[1];
    end
end
assign irqarray5_eventsourceflex81_status = (irqarray5_interrupts[1] | irqarray5_trigger[1]);
always @(*) begin
    irqarray5_eventsourceflex82_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[2]) begin
        if (irqarray5_rising[2]) begin
            irqarray5_eventsourceflex82_trigger_filtered <= (irqarray5_interrupts[2] & (~irqarray5_eventsourceflex82_trigger_d));
        end else begin
            irqarray5_eventsourceflex82_trigger_filtered <= ((~irqarray5_interrupts[2]) & irqarray5_eventsourceflex82_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex82_trigger_filtered <= irqarray5_interrupts[2];
    end
end
assign irqarray5_eventsourceflex82_status = (irqarray5_interrupts[2] | irqarray5_trigger[2]);
always @(*) begin
    irqarray5_eventsourceflex83_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[3]) begin
        if (irqarray5_rising[3]) begin
            irqarray5_eventsourceflex83_trigger_filtered <= (irqarray5_interrupts[3] & (~irqarray5_eventsourceflex83_trigger_d));
        end else begin
            irqarray5_eventsourceflex83_trigger_filtered <= ((~irqarray5_interrupts[3]) & irqarray5_eventsourceflex83_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex83_trigger_filtered <= irqarray5_interrupts[3];
    end
end
assign irqarray5_eventsourceflex83_status = (irqarray5_interrupts[3] | irqarray5_trigger[3]);
always @(*) begin
    irqarray5_eventsourceflex84_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[4]) begin
        if (irqarray5_rising[4]) begin
            irqarray5_eventsourceflex84_trigger_filtered <= (irqarray5_interrupts[4] & (~irqarray5_eventsourceflex84_trigger_d));
        end else begin
            irqarray5_eventsourceflex84_trigger_filtered <= ((~irqarray5_interrupts[4]) & irqarray5_eventsourceflex84_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex84_trigger_filtered <= irqarray5_interrupts[4];
    end
end
assign irqarray5_eventsourceflex84_status = (irqarray5_interrupts[4] | irqarray5_trigger[4]);
always @(*) begin
    irqarray5_eventsourceflex85_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[5]) begin
        if (irqarray5_rising[5]) begin
            irqarray5_eventsourceflex85_trigger_filtered <= (irqarray5_interrupts[5] & (~irqarray5_eventsourceflex85_trigger_d));
        end else begin
            irqarray5_eventsourceflex85_trigger_filtered <= ((~irqarray5_interrupts[5]) & irqarray5_eventsourceflex85_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex85_trigger_filtered <= irqarray5_interrupts[5];
    end
end
assign irqarray5_eventsourceflex85_status = (irqarray5_interrupts[5] | irqarray5_trigger[5]);
always @(*) begin
    irqarray5_eventsourceflex86_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[6]) begin
        if (irqarray5_rising[6]) begin
            irqarray5_eventsourceflex86_trigger_filtered <= (irqarray5_interrupts[6] & (~irqarray5_eventsourceflex86_trigger_d));
        end else begin
            irqarray5_eventsourceflex86_trigger_filtered <= ((~irqarray5_interrupts[6]) & irqarray5_eventsourceflex86_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex86_trigger_filtered <= irqarray5_interrupts[6];
    end
end
assign irqarray5_eventsourceflex86_status = (irqarray5_interrupts[6] | irqarray5_trigger[6]);
always @(*) begin
    irqarray5_eventsourceflex87_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[7]) begin
        if (irqarray5_rising[7]) begin
            irqarray5_eventsourceflex87_trigger_filtered <= (irqarray5_interrupts[7] & (~irqarray5_eventsourceflex87_trigger_d));
        end else begin
            irqarray5_eventsourceflex87_trigger_filtered <= ((~irqarray5_interrupts[7]) & irqarray5_eventsourceflex87_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex87_trigger_filtered <= irqarray5_interrupts[7];
    end
end
assign irqarray5_eventsourceflex87_status = (irqarray5_interrupts[7] | irqarray5_trigger[7]);
always @(*) begin
    irqarray5_eventsourceflex88_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[8]) begin
        if (irqarray5_rising[8]) begin
            irqarray5_eventsourceflex88_trigger_filtered <= (irqarray5_interrupts[8] & (~irqarray5_eventsourceflex88_trigger_d));
        end else begin
            irqarray5_eventsourceflex88_trigger_filtered <= ((~irqarray5_interrupts[8]) & irqarray5_eventsourceflex88_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex88_trigger_filtered <= irqarray5_interrupts[8];
    end
end
assign irqarray5_eventsourceflex88_status = (irqarray5_interrupts[8] | irqarray5_trigger[8]);
always @(*) begin
    irqarray5_eventsourceflex89_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[9]) begin
        if (irqarray5_rising[9]) begin
            irqarray5_eventsourceflex89_trigger_filtered <= (irqarray5_interrupts[9] & (~irqarray5_eventsourceflex89_trigger_d));
        end else begin
            irqarray5_eventsourceflex89_trigger_filtered <= ((~irqarray5_interrupts[9]) & irqarray5_eventsourceflex89_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex89_trigger_filtered <= irqarray5_interrupts[9];
    end
end
assign irqarray5_eventsourceflex89_status = (irqarray5_interrupts[9] | irqarray5_trigger[9]);
always @(*) begin
    irqarray5_eventsourceflex90_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[10]) begin
        if (irqarray5_rising[10]) begin
            irqarray5_eventsourceflex90_trigger_filtered <= (irqarray5_interrupts[10] & (~irqarray5_eventsourceflex90_trigger_d));
        end else begin
            irqarray5_eventsourceflex90_trigger_filtered <= ((~irqarray5_interrupts[10]) & irqarray5_eventsourceflex90_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex90_trigger_filtered <= irqarray5_interrupts[10];
    end
end
assign irqarray5_eventsourceflex90_status = (irqarray5_interrupts[10] | irqarray5_trigger[10]);
always @(*) begin
    irqarray5_eventsourceflex91_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[11]) begin
        if (irqarray5_rising[11]) begin
            irqarray5_eventsourceflex91_trigger_filtered <= (irqarray5_interrupts[11] & (~irqarray5_eventsourceflex91_trigger_d));
        end else begin
            irqarray5_eventsourceflex91_trigger_filtered <= ((~irqarray5_interrupts[11]) & irqarray5_eventsourceflex91_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex91_trigger_filtered <= irqarray5_interrupts[11];
    end
end
assign irqarray5_eventsourceflex91_status = (irqarray5_interrupts[11] | irqarray5_trigger[11]);
always @(*) begin
    irqarray5_eventsourceflex92_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[12]) begin
        if (irqarray5_rising[12]) begin
            irqarray5_eventsourceflex92_trigger_filtered <= (irqarray5_interrupts[12] & (~irqarray5_eventsourceflex92_trigger_d));
        end else begin
            irqarray5_eventsourceflex92_trigger_filtered <= ((~irqarray5_interrupts[12]) & irqarray5_eventsourceflex92_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex92_trigger_filtered <= irqarray5_interrupts[12];
    end
end
assign irqarray5_eventsourceflex92_status = (irqarray5_interrupts[12] | irqarray5_trigger[12]);
always @(*) begin
    irqarray5_eventsourceflex93_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[13]) begin
        if (irqarray5_rising[13]) begin
            irqarray5_eventsourceflex93_trigger_filtered <= (irqarray5_interrupts[13] & (~irqarray5_eventsourceflex93_trigger_d));
        end else begin
            irqarray5_eventsourceflex93_trigger_filtered <= ((~irqarray5_interrupts[13]) & irqarray5_eventsourceflex93_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex93_trigger_filtered <= irqarray5_interrupts[13];
    end
end
assign irqarray5_eventsourceflex93_status = (irqarray5_interrupts[13] | irqarray5_trigger[13]);
always @(*) begin
    irqarray5_eventsourceflex94_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[14]) begin
        if (irqarray5_rising[14]) begin
            irqarray5_eventsourceflex94_trigger_filtered <= (irqarray5_interrupts[14] & (~irqarray5_eventsourceflex94_trigger_d));
        end else begin
            irqarray5_eventsourceflex94_trigger_filtered <= ((~irqarray5_interrupts[14]) & irqarray5_eventsourceflex94_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex94_trigger_filtered <= irqarray5_interrupts[14];
    end
end
assign irqarray5_eventsourceflex94_status = (irqarray5_interrupts[14] | irqarray5_trigger[14]);
always @(*) begin
    irqarray5_eventsourceflex95_trigger_filtered <= 1'd0;
    if (irqarray5_use_edge[15]) begin
        if (irqarray5_rising[15]) begin
            irqarray5_eventsourceflex95_trigger_filtered <= (irqarray5_interrupts[15] & (~irqarray5_eventsourceflex95_trigger_d));
        end else begin
            irqarray5_eventsourceflex95_trigger_filtered <= ((~irqarray5_interrupts[15]) & irqarray5_eventsourceflex95_trigger_d);
        end
    end else begin
        irqarray5_eventsourceflex95_trigger_filtered <= irqarray5_interrupts[15];
    end
end
assign irqarray5_eventsourceflex95_status = (irqarray5_interrupts[15] | irqarray5_trigger[15]);
assign irqarray6_interrupts = irq_remap6;
assign irqarray6_spim0_rx0 = irqarray6_eventsourceflex96_status;
assign irqarray6_spim0_rx1 = irqarray6_eventsourceflex96_pending;
always @(*) begin
    irqarray6_eventsourceflex96_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[0])) begin
        irqarray6_eventsourceflex96_clear <= 1'd1;
    end
end
assign irqarray6_spim0_tx0 = irqarray6_eventsourceflex97_status;
assign irqarray6_spim0_tx1 = irqarray6_eventsourceflex97_pending;
always @(*) begin
    irqarray6_eventsourceflex97_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[1])) begin
        irqarray6_eventsourceflex97_clear <= 1'd1;
    end
end
assign irqarray6_spim0_cmd0 = irqarray6_eventsourceflex98_status;
assign irqarray6_spim0_cmd1 = irqarray6_eventsourceflex98_pending;
always @(*) begin
    irqarray6_eventsourceflex98_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[2])) begin
        irqarray6_eventsourceflex98_clear <= 1'd1;
    end
end
assign irqarray6_spim0_eot0 = irqarray6_eventsourceflex99_status;
assign irqarray6_spim0_eot1 = irqarray6_eventsourceflex99_pending;
always @(*) begin
    irqarray6_eventsourceflex99_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[3])) begin
        irqarray6_eventsourceflex99_clear <= 1'd1;
    end
end
assign irqarray6_spim1_rx0 = irqarray6_eventsourceflex100_status;
assign irqarray6_spim1_rx1 = irqarray6_eventsourceflex100_pending;
always @(*) begin
    irqarray6_eventsourceflex100_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[4])) begin
        irqarray6_eventsourceflex100_clear <= 1'd1;
    end
end
assign irqarray6_spim1_tx0 = irqarray6_eventsourceflex101_status;
assign irqarray6_spim1_tx1 = irqarray6_eventsourceflex101_pending;
always @(*) begin
    irqarray6_eventsourceflex101_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[5])) begin
        irqarray6_eventsourceflex101_clear <= 1'd1;
    end
end
assign irqarray6_spim1_cmd0 = irqarray6_eventsourceflex102_status;
assign irqarray6_spim1_cmd1 = irqarray6_eventsourceflex102_pending;
always @(*) begin
    irqarray6_eventsourceflex102_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[6])) begin
        irqarray6_eventsourceflex102_clear <= 1'd1;
    end
end
assign irqarray6_spim1_eot0 = irqarray6_eventsourceflex103_status;
assign irqarray6_spim1_eot1 = irqarray6_eventsourceflex103_pending;
always @(*) begin
    irqarray6_eventsourceflex103_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[7])) begin
        irqarray6_eventsourceflex103_clear <= 1'd1;
    end
end
assign irqarray6_spim2_rx0 = irqarray6_eventsourceflex104_status;
assign irqarray6_spim2_rx1 = irqarray6_eventsourceflex104_pending;
always @(*) begin
    irqarray6_eventsourceflex104_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[8])) begin
        irqarray6_eventsourceflex104_clear <= 1'd1;
    end
end
assign irqarray6_spim2_tx0 = irqarray6_eventsourceflex105_status;
assign irqarray6_spim2_tx1 = irqarray6_eventsourceflex105_pending;
always @(*) begin
    irqarray6_eventsourceflex105_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[9])) begin
        irqarray6_eventsourceflex105_clear <= 1'd1;
    end
end
assign irqarray6_spim2_cmd0 = irqarray6_eventsourceflex106_status;
assign irqarray6_spim2_cmd1 = irqarray6_eventsourceflex106_pending;
always @(*) begin
    irqarray6_eventsourceflex106_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[10])) begin
        irqarray6_eventsourceflex106_clear <= 1'd1;
    end
end
assign irqarray6_spim2_eot0 = irqarray6_eventsourceflex107_status;
assign irqarray6_spim2_eot1 = irqarray6_eventsourceflex107_pending;
always @(*) begin
    irqarray6_eventsourceflex107_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[11])) begin
        irqarray6_eventsourceflex107_clear <= 1'd1;
    end
end
assign irqarray6_spim3_rx0 = irqarray6_eventsourceflex108_status;
assign irqarray6_spim3_rx1 = irqarray6_eventsourceflex108_pending;
always @(*) begin
    irqarray6_eventsourceflex108_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[12])) begin
        irqarray6_eventsourceflex108_clear <= 1'd1;
    end
end
assign irqarray6_spim3_tx0 = irqarray6_eventsourceflex109_status;
assign irqarray6_spim3_tx1 = irqarray6_eventsourceflex109_pending;
always @(*) begin
    irqarray6_eventsourceflex109_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[13])) begin
        irqarray6_eventsourceflex109_clear <= 1'd1;
    end
end
assign irqarray6_spim3_cmd0 = irqarray6_eventsourceflex110_status;
assign irqarray6_spim3_cmd1 = irqarray6_eventsourceflex110_pending;
always @(*) begin
    irqarray6_eventsourceflex110_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[14])) begin
        irqarray6_eventsourceflex110_clear <= 1'd1;
    end
end
assign irqarray6_spim3_eot0 = irqarray6_eventsourceflex111_status;
assign irqarray6_spim3_eot1 = irqarray6_eventsourceflex111_pending;
always @(*) begin
    irqarray6_eventsourceflex111_clear <= 1'd0;
    if ((irqarray6_pending_re & irqarray6_pending_r[15])) begin
        irqarray6_eventsourceflex111_clear <= 1'd1;
    end
end
assign irqarray6_irq = ((((((((((((((((irqarray6_pending_status[0] & irqarray6_enable_storage[0]) | (irqarray6_pending_status[1] & irqarray6_enable_storage[1])) | (irqarray6_pending_status[2] & irqarray6_enable_storage[2])) | (irqarray6_pending_status[3] & irqarray6_enable_storage[3])) | (irqarray6_pending_status[4] & irqarray6_enable_storage[4])) | (irqarray6_pending_status[5] & irqarray6_enable_storage[5])) | (irqarray6_pending_status[6] & irqarray6_enable_storage[6])) | (irqarray6_pending_status[7] & irqarray6_enable_storage[7])) | (irqarray6_pending_status[8] & irqarray6_enable_storage[8])) | (irqarray6_pending_status[9] & irqarray6_enable_storage[9])) | (irqarray6_pending_status[10] & irqarray6_enable_storage[10])) | (irqarray6_pending_status[11] & irqarray6_enable_storage[11])) | (irqarray6_pending_status[12] & irqarray6_enable_storage[12])) | (irqarray6_pending_status[13] & irqarray6_enable_storage[13])) | (irqarray6_pending_status[14] & irqarray6_enable_storage[14])) | (irqarray6_pending_status[15] & irqarray6_enable_storage[15]));
always @(*) begin
    irqarray6_eventsourceflex96_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[0]) begin
        if (irqarray6_rising[0]) begin
            irqarray6_eventsourceflex96_trigger_filtered <= (irqarray6_interrupts[0] & (~irqarray6_eventsourceflex96_trigger_d));
        end else begin
            irqarray6_eventsourceflex96_trigger_filtered <= ((~irqarray6_interrupts[0]) & irqarray6_eventsourceflex96_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex96_trigger_filtered <= irqarray6_interrupts[0];
    end
end
assign irqarray6_eventsourceflex96_status = (irqarray6_interrupts[0] | irqarray6_trigger[0]);
always @(*) begin
    irqarray6_eventsourceflex97_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[1]) begin
        if (irqarray6_rising[1]) begin
            irqarray6_eventsourceflex97_trigger_filtered <= (irqarray6_interrupts[1] & (~irqarray6_eventsourceflex97_trigger_d));
        end else begin
            irqarray6_eventsourceflex97_trigger_filtered <= ((~irqarray6_interrupts[1]) & irqarray6_eventsourceflex97_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex97_trigger_filtered <= irqarray6_interrupts[1];
    end
end
assign irqarray6_eventsourceflex97_status = (irqarray6_interrupts[1] | irqarray6_trigger[1]);
always @(*) begin
    irqarray6_eventsourceflex98_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[2]) begin
        if (irqarray6_rising[2]) begin
            irqarray6_eventsourceflex98_trigger_filtered <= (irqarray6_interrupts[2] & (~irqarray6_eventsourceflex98_trigger_d));
        end else begin
            irqarray6_eventsourceflex98_trigger_filtered <= ((~irqarray6_interrupts[2]) & irqarray6_eventsourceflex98_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex98_trigger_filtered <= irqarray6_interrupts[2];
    end
end
assign irqarray6_eventsourceflex98_status = (irqarray6_interrupts[2] | irqarray6_trigger[2]);
always @(*) begin
    irqarray6_eventsourceflex99_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[3]) begin
        if (irqarray6_rising[3]) begin
            irqarray6_eventsourceflex99_trigger_filtered <= (irqarray6_interrupts[3] & (~irqarray6_eventsourceflex99_trigger_d));
        end else begin
            irqarray6_eventsourceflex99_trigger_filtered <= ((~irqarray6_interrupts[3]) & irqarray6_eventsourceflex99_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex99_trigger_filtered <= irqarray6_interrupts[3];
    end
end
assign irqarray6_eventsourceflex99_status = (irqarray6_interrupts[3] | irqarray6_trigger[3]);
always @(*) begin
    irqarray6_eventsourceflex100_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[4]) begin
        if (irqarray6_rising[4]) begin
            irqarray6_eventsourceflex100_trigger_filtered <= (irqarray6_interrupts[4] & (~irqarray6_eventsourceflex100_trigger_d));
        end else begin
            irqarray6_eventsourceflex100_trigger_filtered <= ((~irqarray6_interrupts[4]) & irqarray6_eventsourceflex100_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex100_trigger_filtered <= irqarray6_interrupts[4];
    end
end
assign irqarray6_eventsourceflex100_status = (irqarray6_interrupts[4] | irqarray6_trigger[4]);
always @(*) begin
    irqarray6_eventsourceflex101_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[5]) begin
        if (irqarray6_rising[5]) begin
            irqarray6_eventsourceflex101_trigger_filtered <= (irqarray6_interrupts[5] & (~irqarray6_eventsourceflex101_trigger_d));
        end else begin
            irqarray6_eventsourceflex101_trigger_filtered <= ((~irqarray6_interrupts[5]) & irqarray6_eventsourceflex101_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex101_trigger_filtered <= irqarray6_interrupts[5];
    end
end
assign irqarray6_eventsourceflex101_status = (irqarray6_interrupts[5] | irqarray6_trigger[5]);
always @(*) begin
    irqarray6_eventsourceflex102_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[6]) begin
        if (irqarray6_rising[6]) begin
            irqarray6_eventsourceflex102_trigger_filtered <= (irqarray6_interrupts[6] & (~irqarray6_eventsourceflex102_trigger_d));
        end else begin
            irqarray6_eventsourceflex102_trigger_filtered <= ((~irqarray6_interrupts[6]) & irqarray6_eventsourceflex102_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex102_trigger_filtered <= irqarray6_interrupts[6];
    end
end
assign irqarray6_eventsourceflex102_status = (irqarray6_interrupts[6] | irqarray6_trigger[6]);
always @(*) begin
    irqarray6_eventsourceflex103_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[7]) begin
        if (irqarray6_rising[7]) begin
            irqarray6_eventsourceflex103_trigger_filtered <= (irqarray6_interrupts[7] & (~irqarray6_eventsourceflex103_trigger_d));
        end else begin
            irqarray6_eventsourceflex103_trigger_filtered <= ((~irqarray6_interrupts[7]) & irqarray6_eventsourceflex103_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex103_trigger_filtered <= irqarray6_interrupts[7];
    end
end
assign irqarray6_eventsourceflex103_status = (irqarray6_interrupts[7] | irqarray6_trigger[7]);
always @(*) begin
    irqarray6_eventsourceflex104_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[8]) begin
        if (irqarray6_rising[8]) begin
            irqarray6_eventsourceflex104_trigger_filtered <= (irqarray6_interrupts[8] & (~irqarray6_eventsourceflex104_trigger_d));
        end else begin
            irqarray6_eventsourceflex104_trigger_filtered <= ((~irqarray6_interrupts[8]) & irqarray6_eventsourceflex104_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex104_trigger_filtered <= irqarray6_interrupts[8];
    end
end
assign irqarray6_eventsourceflex104_status = (irqarray6_interrupts[8] | irqarray6_trigger[8]);
always @(*) begin
    irqarray6_eventsourceflex105_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[9]) begin
        if (irqarray6_rising[9]) begin
            irqarray6_eventsourceflex105_trigger_filtered <= (irqarray6_interrupts[9] & (~irqarray6_eventsourceflex105_trigger_d));
        end else begin
            irqarray6_eventsourceflex105_trigger_filtered <= ((~irqarray6_interrupts[9]) & irqarray6_eventsourceflex105_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex105_trigger_filtered <= irqarray6_interrupts[9];
    end
end
assign irqarray6_eventsourceflex105_status = (irqarray6_interrupts[9] | irqarray6_trigger[9]);
always @(*) begin
    irqarray6_eventsourceflex106_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[10]) begin
        if (irqarray6_rising[10]) begin
            irqarray6_eventsourceflex106_trigger_filtered <= (irqarray6_interrupts[10] & (~irqarray6_eventsourceflex106_trigger_d));
        end else begin
            irqarray6_eventsourceflex106_trigger_filtered <= ((~irqarray6_interrupts[10]) & irqarray6_eventsourceflex106_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex106_trigger_filtered <= irqarray6_interrupts[10];
    end
end
assign irqarray6_eventsourceflex106_status = (irqarray6_interrupts[10] | irqarray6_trigger[10]);
always @(*) begin
    irqarray6_eventsourceflex107_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[11]) begin
        if (irqarray6_rising[11]) begin
            irqarray6_eventsourceflex107_trigger_filtered <= (irqarray6_interrupts[11] & (~irqarray6_eventsourceflex107_trigger_d));
        end else begin
            irqarray6_eventsourceflex107_trigger_filtered <= ((~irqarray6_interrupts[11]) & irqarray6_eventsourceflex107_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex107_trigger_filtered <= irqarray6_interrupts[11];
    end
end
assign irqarray6_eventsourceflex107_status = (irqarray6_interrupts[11] | irqarray6_trigger[11]);
always @(*) begin
    irqarray6_eventsourceflex108_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[12]) begin
        if (irqarray6_rising[12]) begin
            irqarray6_eventsourceflex108_trigger_filtered <= (irqarray6_interrupts[12] & (~irqarray6_eventsourceflex108_trigger_d));
        end else begin
            irqarray6_eventsourceflex108_trigger_filtered <= ((~irqarray6_interrupts[12]) & irqarray6_eventsourceflex108_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex108_trigger_filtered <= irqarray6_interrupts[12];
    end
end
assign irqarray6_eventsourceflex108_status = (irqarray6_interrupts[12] | irqarray6_trigger[12]);
always @(*) begin
    irqarray6_eventsourceflex109_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[13]) begin
        if (irqarray6_rising[13]) begin
            irqarray6_eventsourceflex109_trigger_filtered <= (irqarray6_interrupts[13] & (~irqarray6_eventsourceflex109_trigger_d));
        end else begin
            irqarray6_eventsourceflex109_trigger_filtered <= ((~irqarray6_interrupts[13]) & irqarray6_eventsourceflex109_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex109_trigger_filtered <= irqarray6_interrupts[13];
    end
end
assign irqarray6_eventsourceflex109_status = (irqarray6_interrupts[13] | irqarray6_trigger[13]);
always @(*) begin
    irqarray6_eventsourceflex110_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[14]) begin
        if (irqarray6_rising[14]) begin
            irqarray6_eventsourceflex110_trigger_filtered <= (irqarray6_interrupts[14] & (~irqarray6_eventsourceflex110_trigger_d));
        end else begin
            irqarray6_eventsourceflex110_trigger_filtered <= ((~irqarray6_interrupts[14]) & irqarray6_eventsourceflex110_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex110_trigger_filtered <= irqarray6_interrupts[14];
    end
end
assign irqarray6_eventsourceflex110_status = (irqarray6_interrupts[14] | irqarray6_trigger[14]);
always @(*) begin
    irqarray6_eventsourceflex111_trigger_filtered <= 1'd0;
    if (irqarray6_use_edge[15]) begin
        if (irqarray6_rising[15]) begin
            irqarray6_eventsourceflex111_trigger_filtered <= (irqarray6_interrupts[15] & (~irqarray6_eventsourceflex111_trigger_d));
        end else begin
            irqarray6_eventsourceflex111_trigger_filtered <= ((~irqarray6_interrupts[15]) & irqarray6_eventsourceflex111_trigger_d);
        end
    end else begin
        irqarray6_eventsourceflex111_trigger_filtered <= irqarray6_interrupts[15];
    end
end
assign irqarray6_eventsourceflex111_status = (irqarray6_interrupts[15] | irqarray6_trigger[15]);
assign irqarray7_interrupts = irq_remap7;
assign irqarray7_i2c0_rx0 = irqarray7_eventsourceflex112_status;
assign irqarray7_i2c0_rx1 = irqarray7_eventsourceflex112_pending;
always @(*) begin
    irqarray7_eventsourceflex112_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[0])) begin
        irqarray7_eventsourceflex112_clear <= 1'd1;
    end
end
assign irqarray7_i2c0_tx0 = irqarray7_eventsourceflex113_status;
assign irqarray7_i2c0_tx1 = irqarray7_eventsourceflex113_pending;
always @(*) begin
    irqarray7_eventsourceflex113_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[1])) begin
        irqarray7_eventsourceflex113_clear <= 1'd1;
    end
end
assign irqarray7_i2c0_cmd0 = irqarray7_eventsourceflex114_status;
assign irqarray7_i2c0_cmd1 = irqarray7_eventsourceflex114_pending;
always @(*) begin
    irqarray7_eventsourceflex114_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[2])) begin
        irqarray7_eventsourceflex114_clear <= 1'd1;
    end
end
assign irqarray7_i2c0_eot0 = irqarray7_eventsourceflex115_status;
assign irqarray7_i2c0_eot1 = irqarray7_eventsourceflex115_pending;
always @(*) begin
    irqarray7_eventsourceflex115_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[3])) begin
        irqarray7_eventsourceflex115_clear <= 1'd1;
    end
end
assign irqarray7_i2c1_rx0 = irqarray7_eventsourceflex116_status;
assign irqarray7_i2c1_rx1 = irqarray7_eventsourceflex116_pending;
always @(*) begin
    irqarray7_eventsourceflex116_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[4])) begin
        irqarray7_eventsourceflex116_clear <= 1'd1;
    end
end
assign irqarray7_i2c1_tx0 = irqarray7_eventsourceflex117_status;
assign irqarray7_i2c1_tx1 = irqarray7_eventsourceflex117_pending;
always @(*) begin
    irqarray7_eventsourceflex117_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[5])) begin
        irqarray7_eventsourceflex117_clear <= 1'd1;
    end
end
assign irqarray7_i2c1_cmd0 = irqarray7_eventsourceflex118_status;
assign irqarray7_i2c1_cmd1 = irqarray7_eventsourceflex118_pending;
always @(*) begin
    irqarray7_eventsourceflex118_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[6])) begin
        irqarray7_eventsourceflex118_clear <= 1'd1;
    end
end
assign irqarray7_i2c1_eot0 = irqarray7_eventsourceflex119_status;
assign irqarray7_i2c1_eot1 = irqarray7_eventsourceflex119_pending;
always @(*) begin
    irqarray7_eventsourceflex119_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[7])) begin
        irqarray7_eventsourceflex119_clear <= 1'd1;
    end
end
assign irqarray7_i2c2_rx0 = irqarray7_eventsourceflex120_status;
assign irqarray7_i2c2_rx1 = irqarray7_eventsourceflex120_pending;
always @(*) begin
    irqarray7_eventsourceflex120_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[8])) begin
        irqarray7_eventsourceflex120_clear <= 1'd1;
    end
end
assign irqarray7_i2c2_tx0 = irqarray7_eventsourceflex121_status;
assign irqarray7_i2c2_tx1 = irqarray7_eventsourceflex121_pending;
always @(*) begin
    irqarray7_eventsourceflex121_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[9])) begin
        irqarray7_eventsourceflex121_clear <= 1'd1;
    end
end
assign irqarray7_i2c2_cmd0 = irqarray7_eventsourceflex122_status;
assign irqarray7_i2c2_cmd1 = irqarray7_eventsourceflex122_pending;
always @(*) begin
    irqarray7_eventsourceflex122_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[10])) begin
        irqarray7_eventsourceflex122_clear <= 1'd1;
    end
end
assign irqarray7_i2c2_eot0 = irqarray7_eventsourceflex123_status;
assign irqarray7_i2c2_eot1 = irqarray7_eventsourceflex123_pending;
always @(*) begin
    irqarray7_eventsourceflex123_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[11])) begin
        irqarray7_eventsourceflex123_clear <= 1'd1;
    end
end
assign irqarray7_i2c3_rx0 = irqarray7_eventsourceflex124_status;
assign irqarray7_i2c3_rx1 = irqarray7_eventsourceflex124_pending;
always @(*) begin
    irqarray7_eventsourceflex124_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[12])) begin
        irqarray7_eventsourceflex124_clear <= 1'd1;
    end
end
assign irqarray7_i2c3_tx0 = irqarray7_eventsourceflex125_status;
assign irqarray7_i2c3_tx1 = irqarray7_eventsourceflex125_pending;
always @(*) begin
    irqarray7_eventsourceflex125_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[13])) begin
        irqarray7_eventsourceflex125_clear <= 1'd1;
    end
end
assign irqarray7_i2c3_cmd0 = irqarray7_eventsourceflex126_status;
assign irqarray7_i2c3_cmd1 = irqarray7_eventsourceflex126_pending;
always @(*) begin
    irqarray7_eventsourceflex126_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[14])) begin
        irqarray7_eventsourceflex126_clear <= 1'd1;
    end
end
assign irqarray7_i2c3_eot0 = irqarray7_eventsourceflex127_status;
assign irqarray7_i2c3_eot1 = irqarray7_eventsourceflex127_pending;
always @(*) begin
    irqarray7_eventsourceflex127_clear <= 1'd0;
    if ((irqarray7_pending_re & irqarray7_pending_r[15])) begin
        irqarray7_eventsourceflex127_clear <= 1'd1;
    end
end
assign irqarray7_irq = ((((((((((((((((irqarray7_pending_status[0] & irqarray7_enable_storage[0]) | (irqarray7_pending_status[1] & irqarray7_enable_storage[1])) | (irqarray7_pending_status[2] & irqarray7_enable_storage[2])) | (irqarray7_pending_status[3] & irqarray7_enable_storage[3])) | (irqarray7_pending_status[4] & irqarray7_enable_storage[4])) | (irqarray7_pending_status[5] & irqarray7_enable_storage[5])) | (irqarray7_pending_status[6] & irqarray7_enable_storage[6])) | (irqarray7_pending_status[7] & irqarray7_enable_storage[7])) | (irqarray7_pending_status[8] & irqarray7_enable_storage[8])) | (irqarray7_pending_status[9] & irqarray7_enable_storage[9])) | (irqarray7_pending_status[10] & irqarray7_enable_storage[10])) | (irqarray7_pending_status[11] & irqarray7_enable_storage[11])) | (irqarray7_pending_status[12] & irqarray7_enable_storage[12])) | (irqarray7_pending_status[13] & irqarray7_enable_storage[13])) | (irqarray7_pending_status[14] & irqarray7_enable_storage[14])) | (irqarray7_pending_status[15] & irqarray7_enable_storage[15]));
always @(*) begin
    irqarray7_eventsourceflex112_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[0]) begin
        if (irqarray7_rising[0]) begin
            irqarray7_eventsourceflex112_trigger_filtered <= (irqarray7_interrupts[0] & (~irqarray7_eventsourceflex112_trigger_d));
        end else begin
            irqarray7_eventsourceflex112_trigger_filtered <= ((~irqarray7_interrupts[0]) & irqarray7_eventsourceflex112_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex112_trigger_filtered <= irqarray7_interrupts[0];
    end
end
assign irqarray7_eventsourceflex112_status = (irqarray7_interrupts[0] | irqarray7_trigger[0]);
always @(*) begin
    irqarray7_eventsourceflex113_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[1]) begin
        if (irqarray7_rising[1]) begin
            irqarray7_eventsourceflex113_trigger_filtered <= (irqarray7_interrupts[1] & (~irqarray7_eventsourceflex113_trigger_d));
        end else begin
            irqarray7_eventsourceflex113_trigger_filtered <= ((~irqarray7_interrupts[1]) & irqarray7_eventsourceflex113_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex113_trigger_filtered <= irqarray7_interrupts[1];
    end
end
assign irqarray7_eventsourceflex113_status = (irqarray7_interrupts[1] | irqarray7_trigger[1]);
always @(*) begin
    irqarray7_eventsourceflex114_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[2]) begin
        if (irqarray7_rising[2]) begin
            irqarray7_eventsourceflex114_trigger_filtered <= (irqarray7_interrupts[2] & (~irqarray7_eventsourceflex114_trigger_d));
        end else begin
            irqarray7_eventsourceflex114_trigger_filtered <= ((~irqarray7_interrupts[2]) & irqarray7_eventsourceflex114_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex114_trigger_filtered <= irqarray7_interrupts[2];
    end
end
assign irqarray7_eventsourceflex114_status = (irqarray7_interrupts[2] | irqarray7_trigger[2]);
always @(*) begin
    irqarray7_eventsourceflex115_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[3]) begin
        if (irqarray7_rising[3]) begin
            irqarray7_eventsourceflex115_trigger_filtered <= (irqarray7_interrupts[3] & (~irqarray7_eventsourceflex115_trigger_d));
        end else begin
            irqarray7_eventsourceflex115_trigger_filtered <= ((~irqarray7_interrupts[3]) & irqarray7_eventsourceflex115_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex115_trigger_filtered <= irqarray7_interrupts[3];
    end
end
assign irqarray7_eventsourceflex115_status = (irqarray7_interrupts[3] | irqarray7_trigger[3]);
always @(*) begin
    irqarray7_eventsourceflex116_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[4]) begin
        if (irqarray7_rising[4]) begin
            irqarray7_eventsourceflex116_trigger_filtered <= (irqarray7_interrupts[4] & (~irqarray7_eventsourceflex116_trigger_d));
        end else begin
            irqarray7_eventsourceflex116_trigger_filtered <= ((~irqarray7_interrupts[4]) & irqarray7_eventsourceflex116_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex116_trigger_filtered <= irqarray7_interrupts[4];
    end
end
assign irqarray7_eventsourceflex116_status = (irqarray7_interrupts[4] | irqarray7_trigger[4]);
always @(*) begin
    irqarray7_eventsourceflex117_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[5]) begin
        if (irqarray7_rising[5]) begin
            irqarray7_eventsourceflex117_trigger_filtered <= (irqarray7_interrupts[5] & (~irqarray7_eventsourceflex117_trigger_d));
        end else begin
            irqarray7_eventsourceflex117_trigger_filtered <= ((~irqarray7_interrupts[5]) & irqarray7_eventsourceflex117_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex117_trigger_filtered <= irqarray7_interrupts[5];
    end
end
assign irqarray7_eventsourceflex117_status = (irqarray7_interrupts[5] | irqarray7_trigger[5]);
always @(*) begin
    irqarray7_eventsourceflex118_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[6]) begin
        if (irqarray7_rising[6]) begin
            irqarray7_eventsourceflex118_trigger_filtered <= (irqarray7_interrupts[6] & (~irqarray7_eventsourceflex118_trigger_d));
        end else begin
            irqarray7_eventsourceflex118_trigger_filtered <= ((~irqarray7_interrupts[6]) & irqarray7_eventsourceflex118_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex118_trigger_filtered <= irqarray7_interrupts[6];
    end
end
assign irqarray7_eventsourceflex118_status = (irqarray7_interrupts[6] | irqarray7_trigger[6]);
always @(*) begin
    irqarray7_eventsourceflex119_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[7]) begin
        if (irqarray7_rising[7]) begin
            irqarray7_eventsourceflex119_trigger_filtered <= (irqarray7_interrupts[7] & (~irqarray7_eventsourceflex119_trigger_d));
        end else begin
            irqarray7_eventsourceflex119_trigger_filtered <= ((~irqarray7_interrupts[7]) & irqarray7_eventsourceflex119_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex119_trigger_filtered <= irqarray7_interrupts[7];
    end
end
assign irqarray7_eventsourceflex119_status = (irqarray7_interrupts[7] | irqarray7_trigger[7]);
always @(*) begin
    irqarray7_eventsourceflex120_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[8]) begin
        if (irqarray7_rising[8]) begin
            irqarray7_eventsourceflex120_trigger_filtered <= (irqarray7_interrupts[8] & (~irqarray7_eventsourceflex120_trigger_d));
        end else begin
            irqarray7_eventsourceflex120_trigger_filtered <= ((~irqarray7_interrupts[8]) & irqarray7_eventsourceflex120_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex120_trigger_filtered <= irqarray7_interrupts[8];
    end
end
assign irqarray7_eventsourceflex120_status = (irqarray7_interrupts[8] | irqarray7_trigger[8]);
always @(*) begin
    irqarray7_eventsourceflex121_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[9]) begin
        if (irqarray7_rising[9]) begin
            irqarray7_eventsourceflex121_trigger_filtered <= (irqarray7_interrupts[9] & (~irqarray7_eventsourceflex121_trigger_d));
        end else begin
            irqarray7_eventsourceflex121_trigger_filtered <= ((~irqarray7_interrupts[9]) & irqarray7_eventsourceflex121_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex121_trigger_filtered <= irqarray7_interrupts[9];
    end
end
assign irqarray7_eventsourceflex121_status = (irqarray7_interrupts[9] | irqarray7_trigger[9]);
always @(*) begin
    irqarray7_eventsourceflex122_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[10]) begin
        if (irqarray7_rising[10]) begin
            irqarray7_eventsourceflex122_trigger_filtered <= (irqarray7_interrupts[10] & (~irqarray7_eventsourceflex122_trigger_d));
        end else begin
            irqarray7_eventsourceflex122_trigger_filtered <= ((~irqarray7_interrupts[10]) & irqarray7_eventsourceflex122_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex122_trigger_filtered <= irqarray7_interrupts[10];
    end
end
assign irqarray7_eventsourceflex122_status = (irqarray7_interrupts[10] | irqarray7_trigger[10]);
always @(*) begin
    irqarray7_eventsourceflex123_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[11]) begin
        if (irqarray7_rising[11]) begin
            irqarray7_eventsourceflex123_trigger_filtered <= (irqarray7_interrupts[11] & (~irqarray7_eventsourceflex123_trigger_d));
        end else begin
            irqarray7_eventsourceflex123_trigger_filtered <= ((~irqarray7_interrupts[11]) & irqarray7_eventsourceflex123_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex123_trigger_filtered <= irqarray7_interrupts[11];
    end
end
assign irqarray7_eventsourceflex123_status = (irqarray7_interrupts[11] | irqarray7_trigger[11]);
always @(*) begin
    irqarray7_eventsourceflex124_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[12]) begin
        if (irqarray7_rising[12]) begin
            irqarray7_eventsourceflex124_trigger_filtered <= (irqarray7_interrupts[12] & (~irqarray7_eventsourceflex124_trigger_d));
        end else begin
            irqarray7_eventsourceflex124_trigger_filtered <= ((~irqarray7_interrupts[12]) & irqarray7_eventsourceflex124_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex124_trigger_filtered <= irqarray7_interrupts[12];
    end
end
assign irqarray7_eventsourceflex124_status = (irqarray7_interrupts[12] | irqarray7_trigger[12]);
always @(*) begin
    irqarray7_eventsourceflex125_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[13]) begin
        if (irqarray7_rising[13]) begin
            irqarray7_eventsourceflex125_trigger_filtered <= (irqarray7_interrupts[13] & (~irqarray7_eventsourceflex125_trigger_d));
        end else begin
            irqarray7_eventsourceflex125_trigger_filtered <= ((~irqarray7_interrupts[13]) & irqarray7_eventsourceflex125_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex125_trigger_filtered <= irqarray7_interrupts[13];
    end
end
assign irqarray7_eventsourceflex125_status = (irqarray7_interrupts[13] | irqarray7_trigger[13]);
always @(*) begin
    irqarray7_eventsourceflex126_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[14]) begin
        if (irqarray7_rising[14]) begin
            irqarray7_eventsourceflex126_trigger_filtered <= (irqarray7_interrupts[14] & (~irqarray7_eventsourceflex126_trigger_d));
        end else begin
            irqarray7_eventsourceflex126_trigger_filtered <= ((~irqarray7_interrupts[14]) & irqarray7_eventsourceflex126_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex126_trigger_filtered <= irqarray7_interrupts[14];
    end
end
assign irqarray7_eventsourceflex126_status = (irqarray7_interrupts[14] | irqarray7_trigger[14]);
always @(*) begin
    irqarray7_eventsourceflex127_trigger_filtered <= 1'd0;
    if (irqarray7_use_edge[15]) begin
        if (irqarray7_rising[15]) begin
            irqarray7_eventsourceflex127_trigger_filtered <= (irqarray7_interrupts[15] & (~irqarray7_eventsourceflex127_trigger_d));
        end else begin
            irqarray7_eventsourceflex127_trigger_filtered <= ((~irqarray7_interrupts[15]) & irqarray7_eventsourceflex127_trigger_d);
        end
    end else begin
        irqarray7_eventsourceflex127_trigger_filtered <= irqarray7_interrupts[15];
    end
end
assign irqarray7_eventsourceflex127_status = (irqarray7_interrupts[15] | irqarray7_trigger[15]);
assign irqarray8_interrupts = irq_remap8;
assign irqarray8_sdio_rx0 = irqarray8_eventsourceflex128_status;
assign irqarray8_sdio_rx1 = irqarray8_eventsourceflex128_pending;
always @(*) begin
    irqarray8_eventsourceflex128_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[0])) begin
        irqarray8_eventsourceflex128_clear <= 1'd1;
    end
end
assign irqarray8_sdio_tx0 = irqarray8_eventsourceflex129_status;
assign irqarray8_sdio_tx1 = irqarray8_eventsourceflex129_pending;
always @(*) begin
    irqarray8_eventsourceflex129_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[1])) begin
        irqarray8_eventsourceflex129_clear <= 1'd1;
    end
end
assign irqarray8_sdio_eot0 = irqarray8_eventsourceflex130_status;
assign irqarray8_sdio_eot1 = irqarray8_eventsourceflex130_pending;
always @(*) begin
    irqarray8_eventsourceflex130_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[2])) begin
        irqarray8_eventsourceflex130_clear <= 1'd1;
    end
end
assign irqarray8_sdio_err0 = irqarray8_eventsourceflex131_status;
assign irqarray8_sdio_err1 = irqarray8_eventsourceflex131_pending;
always @(*) begin
    irqarray8_eventsourceflex131_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[3])) begin
        irqarray8_eventsourceflex131_clear <= 1'd1;
    end
end
assign irqarray8_i2s_rx0 = irqarray8_eventsourceflex132_status;
assign irqarray8_i2s_rx1 = irqarray8_eventsourceflex132_pending;
always @(*) begin
    irqarray8_eventsourceflex132_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[4])) begin
        irqarray8_eventsourceflex132_clear <= 1'd1;
    end
end
assign irqarray8_i2s_tx0 = irqarray8_eventsourceflex133_status;
assign irqarray8_i2s_tx1 = irqarray8_eventsourceflex133_pending;
always @(*) begin
    irqarray8_eventsourceflex133_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[5])) begin
        irqarray8_eventsourceflex133_clear <= 1'd1;
    end
end
assign irqarray8_nc_b8s60 = irqarray8_eventsourceflex134_status;
assign irqarray8_nc_b8s61 = irqarray8_eventsourceflex134_pending;
always @(*) begin
    irqarray8_eventsourceflex134_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[6])) begin
        irqarray8_eventsourceflex134_clear <= 1'd1;
    end
end
assign irqarray8_nc_b8s70 = irqarray8_eventsourceflex135_status;
assign irqarray8_nc_b8s71 = irqarray8_eventsourceflex135_pending;
always @(*) begin
    irqarray8_eventsourceflex135_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[7])) begin
        irqarray8_eventsourceflex135_clear <= 1'd1;
    end
end
assign irqarray8_cam_rx0 = irqarray8_eventsourceflex136_status;
assign irqarray8_cam_rx1 = irqarray8_eventsourceflex136_pending;
always @(*) begin
    irqarray8_eventsourceflex136_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[8])) begin
        irqarray8_eventsourceflex136_clear <= 1'd1;
    end
end
assign irqarray8_adc_rx0 = irqarray8_eventsourceflex137_status;
assign irqarray8_adc_rx1 = irqarray8_eventsourceflex137_pending;
always @(*) begin
    irqarray8_eventsourceflex137_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[9])) begin
        irqarray8_eventsourceflex137_clear <= 1'd1;
    end
end
assign irqarray8_nc_b8s100 = irqarray8_eventsourceflex138_status;
assign irqarray8_nc_b8s101 = irqarray8_eventsourceflex138_pending;
always @(*) begin
    irqarray8_eventsourceflex138_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[10])) begin
        irqarray8_eventsourceflex138_clear <= 1'd1;
    end
end
assign irqarray8_nc_b8s110 = irqarray8_eventsourceflex139_status;
assign irqarray8_nc_b8s111 = irqarray8_eventsourceflex139_pending;
always @(*) begin
    irqarray8_eventsourceflex139_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[11])) begin
        irqarray8_eventsourceflex139_clear <= 1'd1;
    end
end
assign irqarray8_filter_eot0 = irqarray8_eventsourceflex140_status;
assign irqarray8_filter_eot1 = irqarray8_eventsourceflex140_pending;
always @(*) begin
    irqarray8_eventsourceflex140_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[12])) begin
        irqarray8_eventsourceflex140_clear <= 1'd1;
    end
end
assign irqarray8_filter_act0 = irqarray8_eventsourceflex141_status;
assign irqarray8_filter_act1 = irqarray8_eventsourceflex141_pending;
always @(*) begin
    irqarray8_eventsourceflex141_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[13])) begin
        irqarray8_eventsourceflex141_clear <= 1'd1;
    end
end
assign irqarray8_nc_b8s140 = irqarray8_eventsourceflex142_status;
assign irqarray8_nc_b8s141 = irqarray8_eventsourceflex142_pending;
always @(*) begin
    irqarray8_eventsourceflex142_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[14])) begin
        irqarray8_eventsourceflex142_clear <= 1'd1;
    end
end
assign irqarray8_nc_b8s150 = irqarray8_eventsourceflex143_status;
assign irqarray8_nc_b8s151 = irqarray8_eventsourceflex143_pending;
always @(*) begin
    irqarray8_eventsourceflex143_clear <= 1'd0;
    if ((irqarray8_pending_re & irqarray8_pending_r[15])) begin
        irqarray8_eventsourceflex143_clear <= 1'd1;
    end
end
assign irqarray8_irq = ((((((((((((((((irqarray8_pending_status[0] & irqarray8_enable_storage[0]) | (irqarray8_pending_status[1] & irqarray8_enable_storage[1])) | (irqarray8_pending_status[2] & irqarray8_enable_storage[2])) | (irqarray8_pending_status[3] & irqarray8_enable_storage[3])) | (irqarray8_pending_status[4] & irqarray8_enable_storage[4])) | (irqarray8_pending_status[5] & irqarray8_enable_storage[5])) | (irqarray8_pending_status[6] & irqarray8_enable_storage[6])) | (irqarray8_pending_status[7] & irqarray8_enable_storage[7])) | (irqarray8_pending_status[8] & irqarray8_enable_storage[8])) | (irqarray8_pending_status[9] & irqarray8_enable_storage[9])) | (irqarray8_pending_status[10] & irqarray8_enable_storage[10])) | (irqarray8_pending_status[11] & irqarray8_enable_storage[11])) | (irqarray8_pending_status[12] & irqarray8_enable_storage[12])) | (irqarray8_pending_status[13] & irqarray8_enable_storage[13])) | (irqarray8_pending_status[14] & irqarray8_enable_storage[14])) | (irqarray8_pending_status[15] & irqarray8_enable_storage[15]));
always @(*) begin
    irqarray8_eventsourceflex128_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[0]) begin
        if (irqarray8_rising[0]) begin
            irqarray8_eventsourceflex128_trigger_filtered <= (irqarray8_interrupts[0] & (~irqarray8_eventsourceflex128_trigger_d));
        end else begin
            irqarray8_eventsourceflex128_trigger_filtered <= ((~irqarray8_interrupts[0]) & irqarray8_eventsourceflex128_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex128_trigger_filtered <= irqarray8_interrupts[0];
    end
end
assign irqarray8_eventsourceflex128_status = (irqarray8_interrupts[0] | irqarray8_trigger[0]);
always @(*) begin
    irqarray8_eventsourceflex129_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[1]) begin
        if (irqarray8_rising[1]) begin
            irqarray8_eventsourceflex129_trigger_filtered <= (irqarray8_interrupts[1] & (~irqarray8_eventsourceflex129_trigger_d));
        end else begin
            irqarray8_eventsourceflex129_trigger_filtered <= ((~irqarray8_interrupts[1]) & irqarray8_eventsourceflex129_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex129_trigger_filtered <= irqarray8_interrupts[1];
    end
end
assign irqarray8_eventsourceflex129_status = (irqarray8_interrupts[1] | irqarray8_trigger[1]);
always @(*) begin
    irqarray8_eventsourceflex130_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[2]) begin
        if (irqarray8_rising[2]) begin
            irqarray8_eventsourceflex130_trigger_filtered <= (irqarray8_interrupts[2] & (~irqarray8_eventsourceflex130_trigger_d));
        end else begin
            irqarray8_eventsourceflex130_trigger_filtered <= ((~irqarray8_interrupts[2]) & irqarray8_eventsourceflex130_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex130_trigger_filtered <= irqarray8_interrupts[2];
    end
end
assign irqarray8_eventsourceflex130_status = (irqarray8_interrupts[2] | irqarray8_trigger[2]);
always @(*) begin
    irqarray8_eventsourceflex131_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[3]) begin
        if (irqarray8_rising[3]) begin
            irqarray8_eventsourceflex131_trigger_filtered <= (irqarray8_interrupts[3] & (~irqarray8_eventsourceflex131_trigger_d));
        end else begin
            irqarray8_eventsourceflex131_trigger_filtered <= ((~irqarray8_interrupts[3]) & irqarray8_eventsourceflex131_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex131_trigger_filtered <= irqarray8_interrupts[3];
    end
end
assign irqarray8_eventsourceflex131_status = (irqarray8_interrupts[3] | irqarray8_trigger[3]);
always @(*) begin
    irqarray8_eventsourceflex132_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[4]) begin
        if (irqarray8_rising[4]) begin
            irqarray8_eventsourceflex132_trigger_filtered <= (irqarray8_interrupts[4] & (~irqarray8_eventsourceflex132_trigger_d));
        end else begin
            irqarray8_eventsourceflex132_trigger_filtered <= ((~irqarray8_interrupts[4]) & irqarray8_eventsourceflex132_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex132_trigger_filtered <= irqarray8_interrupts[4];
    end
end
assign irqarray8_eventsourceflex132_status = (irqarray8_interrupts[4] | irqarray8_trigger[4]);
always @(*) begin
    irqarray8_eventsourceflex133_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[5]) begin
        if (irqarray8_rising[5]) begin
            irqarray8_eventsourceflex133_trigger_filtered <= (irqarray8_interrupts[5] & (~irqarray8_eventsourceflex133_trigger_d));
        end else begin
            irqarray8_eventsourceflex133_trigger_filtered <= ((~irqarray8_interrupts[5]) & irqarray8_eventsourceflex133_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex133_trigger_filtered <= irqarray8_interrupts[5];
    end
end
assign irqarray8_eventsourceflex133_status = (irqarray8_interrupts[5] | irqarray8_trigger[5]);
always @(*) begin
    irqarray8_eventsourceflex134_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[6]) begin
        if (irqarray8_rising[6]) begin
            irqarray8_eventsourceflex134_trigger_filtered <= (irqarray8_interrupts[6] & (~irqarray8_eventsourceflex134_trigger_d));
        end else begin
            irqarray8_eventsourceflex134_trigger_filtered <= ((~irqarray8_interrupts[6]) & irqarray8_eventsourceflex134_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex134_trigger_filtered <= irqarray8_interrupts[6];
    end
end
assign irqarray8_eventsourceflex134_status = (irqarray8_interrupts[6] | irqarray8_trigger[6]);
always @(*) begin
    irqarray8_eventsourceflex135_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[7]) begin
        if (irqarray8_rising[7]) begin
            irqarray8_eventsourceflex135_trigger_filtered <= (irqarray8_interrupts[7] & (~irqarray8_eventsourceflex135_trigger_d));
        end else begin
            irqarray8_eventsourceflex135_trigger_filtered <= ((~irqarray8_interrupts[7]) & irqarray8_eventsourceflex135_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex135_trigger_filtered <= irqarray8_interrupts[7];
    end
end
assign irqarray8_eventsourceflex135_status = (irqarray8_interrupts[7] | irqarray8_trigger[7]);
always @(*) begin
    irqarray8_eventsourceflex136_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[8]) begin
        if (irqarray8_rising[8]) begin
            irqarray8_eventsourceflex136_trigger_filtered <= (irqarray8_interrupts[8] & (~irqarray8_eventsourceflex136_trigger_d));
        end else begin
            irqarray8_eventsourceflex136_trigger_filtered <= ((~irqarray8_interrupts[8]) & irqarray8_eventsourceflex136_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex136_trigger_filtered <= irqarray8_interrupts[8];
    end
end
assign irqarray8_eventsourceflex136_status = (irqarray8_interrupts[8] | irqarray8_trigger[8]);
always @(*) begin
    irqarray8_eventsourceflex137_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[9]) begin
        if (irqarray8_rising[9]) begin
            irqarray8_eventsourceflex137_trigger_filtered <= (irqarray8_interrupts[9] & (~irqarray8_eventsourceflex137_trigger_d));
        end else begin
            irqarray8_eventsourceflex137_trigger_filtered <= ((~irqarray8_interrupts[9]) & irqarray8_eventsourceflex137_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex137_trigger_filtered <= irqarray8_interrupts[9];
    end
end
assign irqarray8_eventsourceflex137_status = (irqarray8_interrupts[9] | irqarray8_trigger[9]);
always @(*) begin
    irqarray8_eventsourceflex138_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[10]) begin
        if (irqarray8_rising[10]) begin
            irqarray8_eventsourceflex138_trigger_filtered <= (irqarray8_interrupts[10] & (~irqarray8_eventsourceflex138_trigger_d));
        end else begin
            irqarray8_eventsourceflex138_trigger_filtered <= ((~irqarray8_interrupts[10]) & irqarray8_eventsourceflex138_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex138_trigger_filtered <= irqarray8_interrupts[10];
    end
end
assign irqarray8_eventsourceflex138_status = (irqarray8_interrupts[10] | irqarray8_trigger[10]);
always @(*) begin
    irqarray8_eventsourceflex139_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[11]) begin
        if (irqarray8_rising[11]) begin
            irqarray8_eventsourceflex139_trigger_filtered <= (irqarray8_interrupts[11] & (~irqarray8_eventsourceflex139_trigger_d));
        end else begin
            irqarray8_eventsourceflex139_trigger_filtered <= ((~irqarray8_interrupts[11]) & irqarray8_eventsourceflex139_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex139_trigger_filtered <= irqarray8_interrupts[11];
    end
end
assign irqarray8_eventsourceflex139_status = (irqarray8_interrupts[11] | irqarray8_trigger[11]);
always @(*) begin
    irqarray8_eventsourceflex140_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[12]) begin
        if (irqarray8_rising[12]) begin
            irqarray8_eventsourceflex140_trigger_filtered <= (irqarray8_interrupts[12] & (~irqarray8_eventsourceflex140_trigger_d));
        end else begin
            irqarray8_eventsourceflex140_trigger_filtered <= ((~irqarray8_interrupts[12]) & irqarray8_eventsourceflex140_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex140_trigger_filtered <= irqarray8_interrupts[12];
    end
end
assign irqarray8_eventsourceflex140_status = (irqarray8_interrupts[12] | irqarray8_trigger[12]);
always @(*) begin
    irqarray8_eventsourceflex141_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[13]) begin
        if (irqarray8_rising[13]) begin
            irqarray8_eventsourceflex141_trigger_filtered <= (irqarray8_interrupts[13] & (~irqarray8_eventsourceflex141_trigger_d));
        end else begin
            irqarray8_eventsourceflex141_trigger_filtered <= ((~irqarray8_interrupts[13]) & irqarray8_eventsourceflex141_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex141_trigger_filtered <= irqarray8_interrupts[13];
    end
end
assign irqarray8_eventsourceflex141_status = (irqarray8_interrupts[13] | irqarray8_trigger[13]);
always @(*) begin
    irqarray8_eventsourceflex142_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[14]) begin
        if (irqarray8_rising[14]) begin
            irqarray8_eventsourceflex142_trigger_filtered <= (irqarray8_interrupts[14] & (~irqarray8_eventsourceflex142_trigger_d));
        end else begin
            irqarray8_eventsourceflex142_trigger_filtered <= ((~irqarray8_interrupts[14]) & irqarray8_eventsourceflex142_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex142_trigger_filtered <= irqarray8_interrupts[14];
    end
end
assign irqarray8_eventsourceflex142_status = (irqarray8_interrupts[14] | irqarray8_trigger[14]);
always @(*) begin
    irqarray8_eventsourceflex143_trigger_filtered <= 1'd0;
    if (irqarray8_use_edge[15]) begin
        if (irqarray8_rising[15]) begin
            irqarray8_eventsourceflex143_trigger_filtered <= (irqarray8_interrupts[15] & (~irqarray8_eventsourceflex143_trigger_d));
        end else begin
            irqarray8_eventsourceflex143_trigger_filtered <= ((~irqarray8_interrupts[15]) & irqarray8_eventsourceflex143_trigger_d);
        end
    end else begin
        irqarray8_eventsourceflex143_trigger_filtered <= irqarray8_interrupts[15];
    end
end
assign irqarray8_eventsourceflex143_status = (irqarray8_interrupts[15] | irqarray8_trigger[15]);
assign irqarray9_interrupts = irq_remap9;
assign irqarray9_scif_rx0 = irqarray9_eventsourceflex144_status;
assign irqarray9_scif_rx1 = irqarray9_eventsourceflex144_pending;
always @(*) begin
    irqarray9_eventsourceflex144_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[0])) begin
        irqarray9_eventsourceflex144_clear <= 1'd1;
    end
end
assign irqarray9_scif_tx0 = irqarray9_eventsourceflex145_status;
assign irqarray9_scif_tx1 = irqarray9_eventsourceflex145_pending;
always @(*) begin
    irqarray9_eventsourceflex145_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[1])) begin
        irqarray9_eventsourceflex145_clear <= 1'd1;
    end
end
assign irqarray9_scif_rx_char0 = irqarray9_eventsourceflex146_status;
assign irqarray9_scif_rx_char1 = irqarray9_eventsourceflex146_pending;
always @(*) begin
    irqarray9_eventsourceflex146_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[2])) begin
        irqarray9_eventsourceflex146_clear <= 1'd1;
    end
end
assign irqarray9_scif_err0 = irqarray9_eventsourceflex147_status;
assign irqarray9_scif_err1 = irqarray9_eventsourceflex147_pending;
always @(*) begin
    irqarray9_eventsourceflex147_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[3])) begin
        irqarray9_eventsourceflex147_clear <= 1'd1;
    end
end
assign irqarray9_spis0_rx0 = irqarray9_eventsourceflex148_status;
assign irqarray9_spis0_rx1 = irqarray9_eventsourceflex148_pending;
always @(*) begin
    irqarray9_eventsourceflex148_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[4])) begin
        irqarray9_eventsourceflex148_clear <= 1'd1;
    end
end
assign irqarray9_spis0_tx0 = irqarray9_eventsourceflex149_status;
assign irqarray9_spis0_tx1 = irqarray9_eventsourceflex149_pending;
always @(*) begin
    irqarray9_eventsourceflex149_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[5])) begin
        irqarray9_eventsourceflex149_clear <= 1'd1;
    end
end
assign irqarray9_spis0_eot0 = irqarray9_eventsourceflex150_status;
assign irqarray9_spis0_eot1 = irqarray9_eventsourceflex150_pending;
always @(*) begin
    irqarray9_eventsourceflex150_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[6])) begin
        irqarray9_eventsourceflex150_clear <= 1'd1;
    end
end
assign irqarray9_nc_b9s70 = irqarray9_eventsourceflex151_status;
assign irqarray9_nc_b9s71 = irqarray9_eventsourceflex151_pending;
always @(*) begin
    irqarray9_eventsourceflex151_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[7])) begin
        irqarray9_eventsourceflex151_clear <= 1'd1;
    end
end
assign irqarray9_spis1_rx0 = irqarray9_eventsourceflex152_status;
assign irqarray9_spis1_rx1 = irqarray9_eventsourceflex152_pending;
always @(*) begin
    irqarray9_eventsourceflex152_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[8])) begin
        irqarray9_eventsourceflex152_clear <= 1'd1;
    end
end
assign irqarray9_spis1_tx0 = irqarray9_eventsourceflex153_status;
assign irqarray9_spis1_tx1 = irqarray9_eventsourceflex153_pending;
always @(*) begin
    irqarray9_eventsourceflex153_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[9])) begin
        irqarray9_eventsourceflex153_clear <= 1'd1;
    end
end
assign irqarray9_spis1_eot0 = irqarray9_eventsourceflex154_status;
assign irqarray9_spis1_eot1 = irqarray9_eventsourceflex154_pending;
always @(*) begin
    irqarray9_eventsourceflex154_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[10])) begin
        irqarray9_eventsourceflex154_clear <= 1'd1;
    end
end
assign irqarray9_nc_b9s110 = irqarray9_eventsourceflex155_status;
assign irqarray9_nc_b9s111 = irqarray9_eventsourceflex155_pending;
always @(*) begin
    irqarray9_eventsourceflex155_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[11])) begin
        irqarray9_eventsourceflex155_clear <= 1'd1;
    end
end
assign irqarray9_pwm0_ev0 = irqarray9_eventsourceflex156_status;
assign irqarray9_pwm0_ev1 = irqarray9_eventsourceflex156_pending;
always @(*) begin
    irqarray9_eventsourceflex156_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[12])) begin
        irqarray9_eventsourceflex156_clear <= 1'd1;
    end
end
assign irqarray9_pwm1_ev0 = irqarray9_eventsourceflex157_status;
assign irqarray9_pwm1_ev1 = irqarray9_eventsourceflex157_pending;
always @(*) begin
    irqarray9_eventsourceflex157_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[13])) begin
        irqarray9_eventsourceflex157_clear <= 1'd1;
    end
end
assign irqarray9_pwm2_ev0 = irqarray9_eventsourceflex158_status;
assign irqarray9_pwm2_ev1 = irqarray9_eventsourceflex158_pending;
always @(*) begin
    irqarray9_eventsourceflex158_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[14])) begin
        irqarray9_eventsourceflex158_clear <= 1'd1;
    end
end
assign irqarray9_pwm3_ev0 = irqarray9_eventsourceflex159_status;
assign irqarray9_pwm3_ev1 = irqarray9_eventsourceflex159_pending;
always @(*) begin
    irqarray9_eventsourceflex159_clear <= 1'd0;
    if ((irqarray9_pending_re & irqarray9_pending_r[15])) begin
        irqarray9_eventsourceflex159_clear <= 1'd1;
    end
end
assign irqarray9_irq = ((((((((((((((((irqarray9_pending_status[0] & irqarray9_enable_storage[0]) | (irqarray9_pending_status[1] & irqarray9_enable_storage[1])) | (irqarray9_pending_status[2] & irqarray9_enable_storage[2])) | (irqarray9_pending_status[3] & irqarray9_enable_storage[3])) | (irqarray9_pending_status[4] & irqarray9_enable_storage[4])) | (irqarray9_pending_status[5] & irqarray9_enable_storage[5])) | (irqarray9_pending_status[6] & irqarray9_enable_storage[6])) | (irqarray9_pending_status[7] & irqarray9_enable_storage[7])) | (irqarray9_pending_status[8] & irqarray9_enable_storage[8])) | (irqarray9_pending_status[9] & irqarray9_enable_storage[9])) | (irqarray9_pending_status[10] & irqarray9_enable_storage[10])) | (irqarray9_pending_status[11] & irqarray9_enable_storage[11])) | (irqarray9_pending_status[12] & irqarray9_enable_storage[12])) | (irqarray9_pending_status[13] & irqarray9_enable_storage[13])) | (irqarray9_pending_status[14] & irqarray9_enable_storage[14])) | (irqarray9_pending_status[15] & irqarray9_enable_storage[15]));
always @(*) begin
    irqarray9_eventsourceflex144_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[0]) begin
        if (irqarray9_rising[0]) begin
            irqarray9_eventsourceflex144_trigger_filtered <= (irqarray9_interrupts[0] & (~irqarray9_eventsourceflex144_trigger_d));
        end else begin
            irqarray9_eventsourceflex144_trigger_filtered <= ((~irqarray9_interrupts[0]) & irqarray9_eventsourceflex144_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex144_trigger_filtered <= irqarray9_interrupts[0];
    end
end
assign irqarray9_eventsourceflex144_status = (irqarray9_interrupts[0] | irqarray9_trigger[0]);
always @(*) begin
    irqarray9_eventsourceflex145_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[1]) begin
        if (irqarray9_rising[1]) begin
            irqarray9_eventsourceflex145_trigger_filtered <= (irqarray9_interrupts[1] & (~irqarray9_eventsourceflex145_trigger_d));
        end else begin
            irqarray9_eventsourceflex145_trigger_filtered <= ((~irqarray9_interrupts[1]) & irqarray9_eventsourceflex145_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex145_trigger_filtered <= irqarray9_interrupts[1];
    end
end
assign irqarray9_eventsourceflex145_status = (irqarray9_interrupts[1] | irqarray9_trigger[1]);
always @(*) begin
    irqarray9_eventsourceflex146_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[2]) begin
        if (irqarray9_rising[2]) begin
            irqarray9_eventsourceflex146_trigger_filtered <= (irqarray9_interrupts[2] & (~irqarray9_eventsourceflex146_trigger_d));
        end else begin
            irqarray9_eventsourceflex146_trigger_filtered <= ((~irqarray9_interrupts[2]) & irqarray9_eventsourceflex146_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex146_trigger_filtered <= irqarray9_interrupts[2];
    end
end
assign irqarray9_eventsourceflex146_status = (irqarray9_interrupts[2] | irqarray9_trigger[2]);
always @(*) begin
    irqarray9_eventsourceflex147_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[3]) begin
        if (irqarray9_rising[3]) begin
            irqarray9_eventsourceflex147_trigger_filtered <= (irqarray9_interrupts[3] & (~irqarray9_eventsourceflex147_trigger_d));
        end else begin
            irqarray9_eventsourceflex147_trigger_filtered <= ((~irqarray9_interrupts[3]) & irqarray9_eventsourceflex147_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex147_trigger_filtered <= irqarray9_interrupts[3];
    end
end
assign irqarray9_eventsourceflex147_status = (irqarray9_interrupts[3] | irqarray9_trigger[3]);
always @(*) begin
    irqarray9_eventsourceflex148_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[4]) begin
        if (irqarray9_rising[4]) begin
            irqarray9_eventsourceflex148_trigger_filtered <= (irqarray9_interrupts[4] & (~irqarray9_eventsourceflex148_trigger_d));
        end else begin
            irqarray9_eventsourceflex148_trigger_filtered <= ((~irqarray9_interrupts[4]) & irqarray9_eventsourceflex148_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex148_trigger_filtered <= irqarray9_interrupts[4];
    end
end
assign irqarray9_eventsourceflex148_status = (irqarray9_interrupts[4] | irqarray9_trigger[4]);
always @(*) begin
    irqarray9_eventsourceflex149_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[5]) begin
        if (irqarray9_rising[5]) begin
            irqarray9_eventsourceflex149_trigger_filtered <= (irqarray9_interrupts[5] & (~irqarray9_eventsourceflex149_trigger_d));
        end else begin
            irqarray9_eventsourceflex149_trigger_filtered <= ((~irqarray9_interrupts[5]) & irqarray9_eventsourceflex149_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex149_trigger_filtered <= irqarray9_interrupts[5];
    end
end
assign irqarray9_eventsourceflex149_status = (irqarray9_interrupts[5] | irqarray9_trigger[5]);
always @(*) begin
    irqarray9_eventsourceflex150_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[6]) begin
        if (irqarray9_rising[6]) begin
            irqarray9_eventsourceflex150_trigger_filtered <= (irqarray9_interrupts[6] & (~irqarray9_eventsourceflex150_trigger_d));
        end else begin
            irqarray9_eventsourceflex150_trigger_filtered <= ((~irqarray9_interrupts[6]) & irqarray9_eventsourceflex150_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex150_trigger_filtered <= irqarray9_interrupts[6];
    end
end
assign irqarray9_eventsourceflex150_status = (irqarray9_interrupts[6] | irqarray9_trigger[6]);
always @(*) begin
    irqarray9_eventsourceflex151_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[7]) begin
        if (irqarray9_rising[7]) begin
            irqarray9_eventsourceflex151_trigger_filtered <= (irqarray9_interrupts[7] & (~irqarray9_eventsourceflex151_trigger_d));
        end else begin
            irqarray9_eventsourceflex151_trigger_filtered <= ((~irqarray9_interrupts[7]) & irqarray9_eventsourceflex151_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex151_trigger_filtered <= irqarray9_interrupts[7];
    end
end
assign irqarray9_eventsourceflex151_status = (irqarray9_interrupts[7] | irqarray9_trigger[7]);
always @(*) begin
    irqarray9_eventsourceflex152_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[8]) begin
        if (irqarray9_rising[8]) begin
            irqarray9_eventsourceflex152_trigger_filtered <= (irqarray9_interrupts[8] & (~irqarray9_eventsourceflex152_trigger_d));
        end else begin
            irqarray9_eventsourceflex152_trigger_filtered <= ((~irqarray9_interrupts[8]) & irqarray9_eventsourceflex152_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex152_trigger_filtered <= irqarray9_interrupts[8];
    end
end
assign irqarray9_eventsourceflex152_status = (irqarray9_interrupts[8] | irqarray9_trigger[8]);
always @(*) begin
    irqarray9_eventsourceflex153_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[9]) begin
        if (irqarray9_rising[9]) begin
            irqarray9_eventsourceflex153_trigger_filtered <= (irqarray9_interrupts[9] & (~irqarray9_eventsourceflex153_trigger_d));
        end else begin
            irqarray9_eventsourceflex153_trigger_filtered <= ((~irqarray9_interrupts[9]) & irqarray9_eventsourceflex153_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex153_trigger_filtered <= irqarray9_interrupts[9];
    end
end
assign irqarray9_eventsourceflex153_status = (irqarray9_interrupts[9] | irqarray9_trigger[9]);
always @(*) begin
    irqarray9_eventsourceflex154_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[10]) begin
        if (irqarray9_rising[10]) begin
            irqarray9_eventsourceflex154_trigger_filtered <= (irqarray9_interrupts[10] & (~irqarray9_eventsourceflex154_trigger_d));
        end else begin
            irqarray9_eventsourceflex154_trigger_filtered <= ((~irqarray9_interrupts[10]) & irqarray9_eventsourceflex154_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex154_trigger_filtered <= irqarray9_interrupts[10];
    end
end
assign irqarray9_eventsourceflex154_status = (irqarray9_interrupts[10] | irqarray9_trigger[10]);
always @(*) begin
    irqarray9_eventsourceflex155_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[11]) begin
        if (irqarray9_rising[11]) begin
            irqarray9_eventsourceflex155_trigger_filtered <= (irqarray9_interrupts[11] & (~irqarray9_eventsourceflex155_trigger_d));
        end else begin
            irqarray9_eventsourceflex155_trigger_filtered <= ((~irqarray9_interrupts[11]) & irqarray9_eventsourceflex155_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex155_trigger_filtered <= irqarray9_interrupts[11];
    end
end
assign irqarray9_eventsourceflex155_status = (irqarray9_interrupts[11] | irqarray9_trigger[11]);
always @(*) begin
    irqarray9_eventsourceflex156_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[12]) begin
        if (irqarray9_rising[12]) begin
            irqarray9_eventsourceflex156_trigger_filtered <= (irqarray9_interrupts[12] & (~irqarray9_eventsourceflex156_trigger_d));
        end else begin
            irqarray9_eventsourceflex156_trigger_filtered <= ((~irqarray9_interrupts[12]) & irqarray9_eventsourceflex156_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex156_trigger_filtered <= irqarray9_interrupts[12];
    end
end
assign irqarray9_eventsourceflex156_status = (irqarray9_interrupts[12] | irqarray9_trigger[12]);
always @(*) begin
    irqarray9_eventsourceflex157_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[13]) begin
        if (irqarray9_rising[13]) begin
            irqarray9_eventsourceflex157_trigger_filtered <= (irqarray9_interrupts[13] & (~irqarray9_eventsourceflex157_trigger_d));
        end else begin
            irqarray9_eventsourceflex157_trigger_filtered <= ((~irqarray9_interrupts[13]) & irqarray9_eventsourceflex157_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex157_trigger_filtered <= irqarray9_interrupts[13];
    end
end
assign irqarray9_eventsourceflex157_status = (irqarray9_interrupts[13] | irqarray9_trigger[13]);
always @(*) begin
    irqarray9_eventsourceflex158_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[14]) begin
        if (irqarray9_rising[14]) begin
            irqarray9_eventsourceflex158_trigger_filtered <= (irqarray9_interrupts[14] & (~irqarray9_eventsourceflex158_trigger_d));
        end else begin
            irqarray9_eventsourceflex158_trigger_filtered <= ((~irqarray9_interrupts[14]) & irqarray9_eventsourceflex158_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex158_trigger_filtered <= irqarray9_interrupts[14];
    end
end
assign irqarray9_eventsourceflex158_status = (irqarray9_interrupts[14] | irqarray9_trigger[14]);
always @(*) begin
    irqarray9_eventsourceflex159_trigger_filtered <= 1'd0;
    if (irqarray9_use_edge[15]) begin
        if (irqarray9_rising[15]) begin
            irqarray9_eventsourceflex159_trigger_filtered <= (irqarray9_interrupts[15] & (~irqarray9_eventsourceflex159_trigger_d));
        end else begin
            irqarray9_eventsourceflex159_trigger_filtered <= ((~irqarray9_interrupts[15]) & irqarray9_eventsourceflex159_trigger_d);
        end
    end else begin
        irqarray9_eventsourceflex159_trigger_filtered <= irqarray9_interrupts[15];
    end
end
assign irqarray9_eventsourceflex159_status = (irqarray9_interrupts[15] | irqarray9_trigger[15]);
assign irqarray10_interrupts = irq_remap10;
assign irqarray10_ioxirq0 = irqarray10_eventsourceflex160_status;
assign irqarray10_ioxirq1 = irqarray10_eventsourceflex160_pending;
always @(*) begin
    irqarray10_eventsourceflex160_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[0])) begin
        irqarray10_eventsourceflex160_clear <= 1'd1;
    end
end
assign irqarray10_usbc0 = irqarray10_eventsourceflex161_status;
assign irqarray10_usbc1 = irqarray10_eventsourceflex161_pending;
always @(*) begin
    irqarray10_eventsourceflex161_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[1])) begin
        irqarray10_eventsourceflex161_clear <= 1'd1;
    end
end
assign irqarray10_sddcirq0 = irqarray10_eventsourceflex162_status;
assign irqarray10_sddcirq1 = irqarray10_eventsourceflex162_pending;
always @(*) begin
    irqarray10_eventsourceflex162_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[2])) begin
        irqarray10_eventsourceflex162_clear <= 1'd1;
    end
end
assign irqarray10_pioirq00 = irqarray10_eventsourceflex163_status;
assign irqarray10_pioirq01 = irqarray10_eventsourceflex163_pending;
always @(*) begin
    irqarray10_eventsourceflex163_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[3])) begin
        irqarray10_eventsourceflex163_clear <= 1'd1;
    end
end
assign irqarray10_pioirq10 = irqarray10_eventsourceflex164_status;
assign irqarray10_pioirq11 = irqarray10_eventsourceflex164_pending;
always @(*) begin
    irqarray10_eventsourceflex164_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[4])) begin
        irqarray10_eventsourceflex164_clear <= 1'd1;
    end
end
assign irqarray10_pioirq20 = irqarray10_eventsourceflex165_status;
assign irqarray10_pioirq21 = irqarray10_eventsourceflex165_pending;
always @(*) begin
    irqarray10_eventsourceflex165_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[5])) begin
        irqarray10_eventsourceflex165_clear <= 1'd1;
    end
end
assign irqarray10_pioirq30 = irqarray10_eventsourceflex166_status;
assign irqarray10_pioirq31 = irqarray10_eventsourceflex166_pending;
always @(*) begin
    irqarray10_eventsourceflex166_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[6])) begin
        irqarray10_eventsourceflex166_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s70 = irqarray10_eventsourceflex167_status;
assign irqarray10_nc_b10s71 = irqarray10_eventsourceflex167_pending;
always @(*) begin
    irqarray10_eventsourceflex167_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[7])) begin
        irqarray10_eventsourceflex167_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s80 = irqarray10_eventsourceflex168_status;
assign irqarray10_nc_b10s81 = irqarray10_eventsourceflex168_pending;
always @(*) begin
    irqarray10_eventsourceflex168_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[8])) begin
        irqarray10_eventsourceflex168_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s90 = irqarray10_eventsourceflex169_status;
assign irqarray10_nc_b10s91 = irqarray10_eventsourceflex169_pending;
always @(*) begin
    irqarray10_eventsourceflex169_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[9])) begin
        irqarray10_eventsourceflex169_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s100 = irqarray10_eventsourceflex170_status;
assign irqarray10_nc_b10s101 = irqarray10_eventsourceflex170_pending;
always @(*) begin
    irqarray10_eventsourceflex170_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[10])) begin
        irqarray10_eventsourceflex170_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s110 = irqarray10_eventsourceflex171_status;
assign irqarray10_nc_b10s111 = irqarray10_eventsourceflex171_pending;
always @(*) begin
    irqarray10_eventsourceflex171_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[11])) begin
        irqarray10_eventsourceflex171_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s120 = irqarray10_eventsourceflex172_status;
assign irqarray10_nc_b10s121 = irqarray10_eventsourceflex172_pending;
always @(*) begin
    irqarray10_eventsourceflex172_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[12])) begin
        irqarray10_eventsourceflex172_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s130 = irqarray10_eventsourceflex173_status;
assign irqarray10_nc_b10s131 = irqarray10_eventsourceflex173_pending;
always @(*) begin
    irqarray10_eventsourceflex173_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[13])) begin
        irqarray10_eventsourceflex173_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s140 = irqarray10_eventsourceflex174_status;
assign irqarray10_nc_b10s141 = irqarray10_eventsourceflex174_pending;
always @(*) begin
    irqarray10_eventsourceflex174_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[14])) begin
        irqarray10_eventsourceflex174_clear <= 1'd1;
    end
end
assign irqarray10_nc_b10s150 = irqarray10_eventsourceflex175_status;
assign irqarray10_nc_b10s151 = irqarray10_eventsourceflex175_pending;
always @(*) begin
    irqarray10_eventsourceflex175_clear <= 1'd0;
    if ((irqarray10_pending_re & irqarray10_pending_r[15])) begin
        irqarray10_eventsourceflex175_clear <= 1'd1;
    end
end
assign irqarray10_irq = ((((((((((((((((irqarray10_pending_status[0] & irqarray10_enable_storage[0]) | (irqarray10_pending_status[1] & irqarray10_enable_storage[1])) | (irqarray10_pending_status[2] & irqarray10_enable_storage[2])) | (irqarray10_pending_status[3] & irqarray10_enable_storage[3])) | (irqarray10_pending_status[4] & irqarray10_enable_storage[4])) | (irqarray10_pending_status[5] & irqarray10_enable_storage[5])) | (irqarray10_pending_status[6] & irqarray10_enable_storage[6])) | (irqarray10_pending_status[7] & irqarray10_enable_storage[7])) | (irqarray10_pending_status[8] & irqarray10_enable_storage[8])) | (irqarray10_pending_status[9] & irqarray10_enable_storage[9])) | (irqarray10_pending_status[10] & irqarray10_enable_storage[10])) | (irqarray10_pending_status[11] & irqarray10_enable_storage[11])) | (irqarray10_pending_status[12] & irqarray10_enable_storage[12])) | (irqarray10_pending_status[13] & irqarray10_enable_storage[13])) | (irqarray10_pending_status[14] & irqarray10_enable_storage[14])) | (irqarray10_pending_status[15] & irqarray10_enable_storage[15]));
always @(*) begin
    irqarray10_eventsourceflex160_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[0]) begin
        if (irqarray10_rising[0]) begin
            irqarray10_eventsourceflex160_trigger_filtered <= (irqarray10_interrupts[0] & (~irqarray10_eventsourceflex160_trigger_d));
        end else begin
            irqarray10_eventsourceflex160_trigger_filtered <= ((~irqarray10_interrupts[0]) & irqarray10_eventsourceflex160_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex160_trigger_filtered <= irqarray10_interrupts[0];
    end
end
assign irqarray10_eventsourceflex160_status = (irqarray10_interrupts[0] | irqarray10_trigger[0]);
always @(*) begin
    irqarray10_eventsourceflex161_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[1]) begin
        if (irqarray10_rising[1]) begin
            irqarray10_eventsourceflex161_trigger_filtered <= (irqarray10_interrupts[1] & (~irqarray10_eventsourceflex161_trigger_d));
        end else begin
            irqarray10_eventsourceflex161_trigger_filtered <= ((~irqarray10_interrupts[1]) & irqarray10_eventsourceflex161_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex161_trigger_filtered <= irqarray10_interrupts[1];
    end
end
assign irqarray10_eventsourceflex161_status = (irqarray10_interrupts[1] | irqarray10_trigger[1]);
always @(*) begin
    irqarray10_eventsourceflex162_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[2]) begin
        if (irqarray10_rising[2]) begin
            irqarray10_eventsourceflex162_trigger_filtered <= (irqarray10_interrupts[2] & (~irqarray10_eventsourceflex162_trigger_d));
        end else begin
            irqarray10_eventsourceflex162_trigger_filtered <= ((~irqarray10_interrupts[2]) & irqarray10_eventsourceflex162_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex162_trigger_filtered <= irqarray10_interrupts[2];
    end
end
assign irqarray10_eventsourceflex162_status = (irqarray10_interrupts[2] | irqarray10_trigger[2]);
always @(*) begin
    irqarray10_eventsourceflex163_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[3]) begin
        if (irqarray10_rising[3]) begin
            irqarray10_eventsourceflex163_trigger_filtered <= (irqarray10_interrupts[3] & (~irqarray10_eventsourceflex163_trigger_d));
        end else begin
            irqarray10_eventsourceflex163_trigger_filtered <= ((~irqarray10_interrupts[3]) & irqarray10_eventsourceflex163_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex163_trigger_filtered <= irqarray10_interrupts[3];
    end
end
assign irqarray10_eventsourceflex163_status = (irqarray10_interrupts[3] | irqarray10_trigger[3]);
always @(*) begin
    irqarray10_eventsourceflex164_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[4]) begin
        if (irqarray10_rising[4]) begin
            irqarray10_eventsourceflex164_trigger_filtered <= (irqarray10_interrupts[4] & (~irqarray10_eventsourceflex164_trigger_d));
        end else begin
            irqarray10_eventsourceflex164_trigger_filtered <= ((~irqarray10_interrupts[4]) & irqarray10_eventsourceflex164_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex164_trigger_filtered <= irqarray10_interrupts[4];
    end
end
assign irqarray10_eventsourceflex164_status = (irqarray10_interrupts[4] | irqarray10_trigger[4]);
always @(*) begin
    irqarray10_eventsourceflex165_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[5]) begin
        if (irqarray10_rising[5]) begin
            irqarray10_eventsourceflex165_trigger_filtered <= (irqarray10_interrupts[5] & (~irqarray10_eventsourceflex165_trigger_d));
        end else begin
            irqarray10_eventsourceflex165_trigger_filtered <= ((~irqarray10_interrupts[5]) & irqarray10_eventsourceflex165_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex165_trigger_filtered <= irqarray10_interrupts[5];
    end
end
assign irqarray10_eventsourceflex165_status = (irqarray10_interrupts[5] | irqarray10_trigger[5]);
always @(*) begin
    irqarray10_eventsourceflex166_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[6]) begin
        if (irqarray10_rising[6]) begin
            irqarray10_eventsourceflex166_trigger_filtered <= (irqarray10_interrupts[6] & (~irqarray10_eventsourceflex166_trigger_d));
        end else begin
            irqarray10_eventsourceflex166_trigger_filtered <= ((~irqarray10_interrupts[6]) & irqarray10_eventsourceflex166_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex166_trigger_filtered <= irqarray10_interrupts[6];
    end
end
assign irqarray10_eventsourceflex166_status = (irqarray10_interrupts[6] | irqarray10_trigger[6]);
always @(*) begin
    irqarray10_eventsourceflex167_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[7]) begin
        if (irqarray10_rising[7]) begin
            irqarray10_eventsourceflex167_trigger_filtered <= (irqarray10_interrupts[7] & (~irqarray10_eventsourceflex167_trigger_d));
        end else begin
            irqarray10_eventsourceflex167_trigger_filtered <= ((~irqarray10_interrupts[7]) & irqarray10_eventsourceflex167_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex167_trigger_filtered <= irqarray10_interrupts[7];
    end
end
assign irqarray10_eventsourceflex167_status = (irqarray10_interrupts[7] | irqarray10_trigger[7]);
always @(*) begin
    irqarray10_eventsourceflex168_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[8]) begin
        if (irqarray10_rising[8]) begin
            irqarray10_eventsourceflex168_trigger_filtered <= (irqarray10_interrupts[8] & (~irqarray10_eventsourceflex168_trigger_d));
        end else begin
            irqarray10_eventsourceflex168_trigger_filtered <= ((~irqarray10_interrupts[8]) & irqarray10_eventsourceflex168_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex168_trigger_filtered <= irqarray10_interrupts[8];
    end
end
assign irqarray10_eventsourceflex168_status = (irqarray10_interrupts[8] | irqarray10_trigger[8]);
always @(*) begin
    irqarray10_eventsourceflex169_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[9]) begin
        if (irqarray10_rising[9]) begin
            irqarray10_eventsourceflex169_trigger_filtered <= (irqarray10_interrupts[9] & (~irqarray10_eventsourceflex169_trigger_d));
        end else begin
            irqarray10_eventsourceflex169_trigger_filtered <= ((~irqarray10_interrupts[9]) & irqarray10_eventsourceflex169_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex169_trigger_filtered <= irqarray10_interrupts[9];
    end
end
assign irqarray10_eventsourceflex169_status = (irqarray10_interrupts[9] | irqarray10_trigger[9]);
always @(*) begin
    irqarray10_eventsourceflex170_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[10]) begin
        if (irqarray10_rising[10]) begin
            irqarray10_eventsourceflex170_trigger_filtered <= (irqarray10_interrupts[10] & (~irqarray10_eventsourceflex170_trigger_d));
        end else begin
            irqarray10_eventsourceflex170_trigger_filtered <= ((~irqarray10_interrupts[10]) & irqarray10_eventsourceflex170_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex170_trigger_filtered <= irqarray10_interrupts[10];
    end
end
assign irqarray10_eventsourceflex170_status = (irqarray10_interrupts[10] | irqarray10_trigger[10]);
always @(*) begin
    irqarray10_eventsourceflex171_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[11]) begin
        if (irqarray10_rising[11]) begin
            irqarray10_eventsourceflex171_trigger_filtered <= (irqarray10_interrupts[11] & (~irqarray10_eventsourceflex171_trigger_d));
        end else begin
            irqarray10_eventsourceflex171_trigger_filtered <= ((~irqarray10_interrupts[11]) & irqarray10_eventsourceflex171_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex171_trigger_filtered <= irqarray10_interrupts[11];
    end
end
assign irqarray10_eventsourceflex171_status = (irqarray10_interrupts[11] | irqarray10_trigger[11]);
always @(*) begin
    irqarray10_eventsourceflex172_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[12]) begin
        if (irqarray10_rising[12]) begin
            irqarray10_eventsourceflex172_trigger_filtered <= (irqarray10_interrupts[12] & (~irqarray10_eventsourceflex172_trigger_d));
        end else begin
            irqarray10_eventsourceflex172_trigger_filtered <= ((~irqarray10_interrupts[12]) & irqarray10_eventsourceflex172_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex172_trigger_filtered <= irqarray10_interrupts[12];
    end
end
assign irqarray10_eventsourceflex172_status = (irqarray10_interrupts[12] | irqarray10_trigger[12]);
always @(*) begin
    irqarray10_eventsourceflex173_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[13]) begin
        if (irqarray10_rising[13]) begin
            irqarray10_eventsourceflex173_trigger_filtered <= (irqarray10_interrupts[13] & (~irqarray10_eventsourceflex173_trigger_d));
        end else begin
            irqarray10_eventsourceflex173_trigger_filtered <= ((~irqarray10_interrupts[13]) & irqarray10_eventsourceflex173_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex173_trigger_filtered <= irqarray10_interrupts[13];
    end
end
assign irqarray10_eventsourceflex173_status = (irqarray10_interrupts[13] | irqarray10_trigger[13]);
always @(*) begin
    irqarray10_eventsourceflex174_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[14]) begin
        if (irqarray10_rising[14]) begin
            irqarray10_eventsourceflex174_trigger_filtered <= (irqarray10_interrupts[14] & (~irqarray10_eventsourceflex174_trigger_d));
        end else begin
            irqarray10_eventsourceflex174_trigger_filtered <= ((~irqarray10_interrupts[14]) & irqarray10_eventsourceflex174_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex174_trigger_filtered <= irqarray10_interrupts[14];
    end
end
assign irqarray10_eventsourceflex174_status = (irqarray10_interrupts[14] | irqarray10_trigger[14]);
always @(*) begin
    irqarray10_eventsourceflex175_trigger_filtered <= 1'd0;
    if (irqarray10_use_edge[15]) begin
        if (irqarray10_rising[15]) begin
            irqarray10_eventsourceflex175_trigger_filtered <= (irqarray10_interrupts[15] & (~irqarray10_eventsourceflex175_trigger_d));
        end else begin
            irqarray10_eventsourceflex175_trigger_filtered <= ((~irqarray10_interrupts[15]) & irqarray10_eventsourceflex175_trigger_d);
        end
    end else begin
        irqarray10_eventsourceflex175_trigger_filtered <= irqarray10_interrupts[15];
    end
end
assign irqarray10_eventsourceflex175_status = (irqarray10_interrupts[15] | irqarray10_trigger[15]);
assign irqarray11_interrupts = irq_remap11;
assign irqarray11_i2s_rx_dupe0 = irqarray11_eventsourceflex176_status;
assign irqarray11_i2s_rx_dupe1 = irqarray11_eventsourceflex176_pending;
always @(*) begin
    irqarray11_eventsourceflex176_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[0])) begin
        irqarray11_eventsourceflex176_clear <= 1'd1;
    end
end
assign irqarray11_i2s_tx_dupe0 = irqarray11_eventsourceflex177_status;
assign irqarray11_i2s_tx_dupe1 = irqarray11_eventsourceflex177_pending;
always @(*) begin
    irqarray11_eventsourceflex177_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[1])) begin
        irqarray11_eventsourceflex177_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s20 = irqarray11_eventsourceflex178_status;
assign irqarray11_nc_b11s21 = irqarray11_eventsourceflex178_pending;
always @(*) begin
    irqarray11_eventsourceflex178_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[2])) begin
        irqarray11_eventsourceflex178_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s30 = irqarray11_eventsourceflex179_status;
assign irqarray11_nc_b11s31 = irqarray11_eventsourceflex179_pending;
always @(*) begin
    irqarray11_eventsourceflex179_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[3])) begin
        irqarray11_eventsourceflex179_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s40 = irqarray11_eventsourceflex180_status;
assign irqarray11_nc_b11s41 = irqarray11_eventsourceflex180_pending;
always @(*) begin
    irqarray11_eventsourceflex180_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[4])) begin
        irqarray11_eventsourceflex180_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s50 = irqarray11_eventsourceflex181_status;
assign irqarray11_nc_b11s51 = irqarray11_eventsourceflex181_pending;
always @(*) begin
    irqarray11_eventsourceflex181_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[5])) begin
        irqarray11_eventsourceflex181_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s60 = irqarray11_eventsourceflex182_status;
assign irqarray11_nc_b11s61 = irqarray11_eventsourceflex182_pending;
always @(*) begin
    irqarray11_eventsourceflex182_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[6])) begin
        irqarray11_eventsourceflex182_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s70 = irqarray11_eventsourceflex183_status;
assign irqarray11_nc_b11s71 = irqarray11_eventsourceflex183_pending;
always @(*) begin
    irqarray11_eventsourceflex183_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[7])) begin
        irqarray11_eventsourceflex183_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s80 = irqarray11_eventsourceflex184_status;
assign irqarray11_nc_b11s81 = irqarray11_eventsourceflex184_pending;
always @(*) begin
    irqarray11_eventsourceflex184_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[8])) begin
        irqarray11_eventsourceflex184_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s90 = irqarray11_eventsourceflex185_status;
assign irqarray11_nc_b11s91 = irqarray11_eventsourceflex185_pending;
always @(*) begin
    irqarray11_eventsourceflex185_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[9])) begin
        irqarray11_eventsourceflex185_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s100 = irqarray11_eventsourceflex186_status;
assign irqarray11_nc_b11s101 = irqarray11_eventsourceflex186_pending;
always @(*) begin
    irqarray11_eventsourceflex186_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[10])) begin
        irqarray11_eventsourceflex186_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s110 = irqarray11_eventsourceflex187_status;
assign irqarray11_nc_b11s111 = irqarray11_eventsourceflex187_pending;
always @(*) begin
    irqarray11_eventsourceflex187_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[11])) begin
        irqarray11_eventsourceflex187_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s120 = irqarray11_eventsourceflex188_status;
assign irqarray11_nc_b11s121 = irqarray11_eventsourceflex188_pending;
always @(*) begin
    irqarray11_eventsourceflex188_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[12])) begin
        irqarray11_eventsourceflex188_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s130 = irqarray11_eventsourceflex189_status;
assign irqarray11_nc_b11s131 = irqarray11_eventsourceflex189_pending;
always @(*) begin
    irqarray11_eventsourceflex189_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[13])) begin
        irqarray11_eventsourceflex189_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s140 = irqarray11_eventsourceflex190_status;
assign irqarray11_nc_b11s141 = irqarray11_eventsourceflex190_pending;
always @(*) begin
    irqarray11_eventsourceflex190_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[14])) begin
        irqarray11_eventsourceflex190_clear <= 1'd1;
    end
end
assign irqarray11_nc_b11s150 = irqarray11_eventsourceflex191_status;
assign irqarray11_nc_b11s151 = irqarray11_eventsourceflex191_pending;
always @(*) begin
    irqarray11_eventsourceflex191_clear <= 1'd0;
    if ((irqarray11_pending_re & irqarray11_pending_r[15])) begin
        irqarray11_eventsourceflex191_clear <= 1'd1;
    end
end
assign irqarray11_irq = ((((((((((((((((irqarray11_pending_status[0] & irqarray11_enable_storage[0]) | (irqarray11_pending_status[1] & irqarray11_enable_storage[1])) | (irqarray11_pending_status[2] & irqarray11_enable_storage[2])) | (irqarray11_pending_status[3] & irqarray11_enable_storage[3])) | (irqarray11_pending_status[4] & irqarray11_enable_storage[4])) | (irqarray11_pending_status[5] & irqarray11_enable_storage[5])) | (irqarray11_pending_status[6] & irqarray11_enable_storage[6])) | (irqarray11_pending_status[7] & irqarray11_enable_storage[7])) | (irqarray11_pending_status[8] & irqarray11_enable_storage[8])) | (irqarray11_pending_status[9] & irqarray11_enable_storage[9])) | (irqarray11_pending_status[10] & irqarray11_enable_storage[10])) | (irqarray11_pending_status[11] & irqarray11_enable_storage[11])) | (irqarray11_pending_status[12] & irqarray11_enable_storage[12])) | (irqarray11_pending_status[13] & irqarray11_enable_storage[13])) | (irqarray11_pending_status[14] & irqarray11_enable_storage[14])) | (irqarray11_pending_status[15] & irqarray11_enable_storage[15]));
always @(*) begin
    irqarray11_eventsourceflex176_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[0]) begin
        if (irqarray11_rising[0]) begin
            irqarray11_eventsourceflex176_trigger_filtered <= (irqarray11_interrupts[0] & (~irqarray11_eventsourceflex176_trigger_d));
        end else begin
            irqarray11_eventsourceflex176_trigger_filtered <= ((~irqarray11_interrupts[0]) & irqarray11_eventsourceflex176_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex176_trigger_filtered <= irqarray11_interrupts[0];
    end
end
assign irqarray11_eventsourceflex176_status = (irqarray11_interrupts[0] | irqarray11_trigger[0]);
always @(*) begin
    irqarray11_eventsourceflex177_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[1]) begin
        if (irqarray11_rising[1]) begin
            irqarray11_eventsourceflex177_trigger_filtered <= (irqarray11_interrupts[1] & (~irqarray11_eventsourceflex177_trigger_d));
        end else begin
            irqarray11_eventsourceflex177_trigger_filtered <= ((~irqarray11_interrupts[1]) & irqarray11_eventsourceflex177_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex177_trigger_filtered <= irqarray11_interrupts[1];
    end
end
assign irqarray11_eventsourceflex177_status = (irqarray11_interrupts[1] | irqarray11_trigger[1]);
always @(*) begin
    irqarray11_eventsourceflex178_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[2]) begin
        if (irqarray11_rising[2]) begin
            irqarray11_eventsourceflex178_trigger_filtered <= (irqarray11_interrupts[2] & (~irqarray11_eventsourceflex178_trigger_d));
        end else begin
            irqarray11_eventsourceflex178_trigger_filtered <= ((~irqarray11_interrupts[2]) & irqarray11_eventsourceflex178_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex178_trigger_filtered <= irqarray11_interrupts[2];
    end
end
assign irqarray11_eventsourceflex178_status = (irqarray11_interrupts[2] | irqarray11_trigger[2]);
always @(*) begin
    irqarray11_eventsourceflex179_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[3]) begin
        if (irqarray11_rising[3]) begin
            irqarray11_eventsourceflex179_trigger_filtered <= (irqarray11_interrupts[3] & (~irqarray11_eventsourceflex179_trigger_d));
        end else begin
            irqarray11_eventsourceflex179_trigger_filtered <= ((~irqarray11_interrupts[3]) & irqarray11_eventsourceflex179_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex179_trigger_filtered <= irqarray11_interrupts[3];
    end
end
assign irqarray11_eventsourceflex179_status = (irqarray11_interrupts[3] | irqarray11_trigger[3]);
always @(*) begin
    irqarray11_eventsourceflex180_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[4]) begin
        if (irqarray11_rising[4]) begin
            irqarray11_eventsourceflex180_trigger_filtered <= (irqarray11_interrupts[4] & (~irqarray11_eventsourceflex180_trigger_d));
        end else begin
            irqarray11_eventsourceflex180_trigger_filtered <= ((~irqarray11_interrupts[4]) & irqarray11_eventsourceflex180_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex180_trigger_filtered <= irqarray11_interrupts[4];
    end
end
assign irqarray11_eventsourceflex180_status = (irqarray11_interrupts[4] | irqarray11_trigger[4]);
always @(*) begin
    irqarray11_eventsourceflex181_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[5]) begin
        if (irqarray11_rising[5]) begin
            irqarray11_eventsourceflex181_trigger_filtered <= (irqarray11_interrupts[5] & (~irqarray11_eventsourceflex181_trigger_d));
        end else begin
            irqarray11_eventsourceflex181_trigger_filtered <= ((~irqarray11_interrupts[5]) & irqarray11_eventsourceflex181_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex181_trigger_filtered <= irqarray11_interrupts[5];
    end
end
assign irqarray11_eventsourceflex181_status = (irqarray11_interrupts[5] | irqarray11_trigger[5]);
always @(*) begin
    irqarray11_eventsourceflex182_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[6]) begin
        if (irqarray11_rising[6]) begin
            irqarray11_eventsourceflex182_trigger_filtered <= (irqarray11_interrupts[6] & (~irqarray11_eventsourceflex182_trigger_d));
        end else begin
            irqarray11_eventsourceflex182_trigger_filtered <= ((~irqarray11_interrupts[6]) & irqarray11_eventsourceflex182_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex182_trigger_filtered <= irqarray11_interrupts[6];
    end
end
assign irqarray11_eventsourceflex182_status = (irqarray11_interrupts[6] | irqarray11_trigger[6]);
always @(*) begin
    irqarray11_eventsourceflex183_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[7]) begin
        if (irqarray11_rising[7]) begin
            irqarray11_eventsourceflex183_trigger_filtered <= (irqarray11_interrupts[7] & (~irqarray11_eventsourceflex183_trigger_d));
        end else begin
            irqarray11_eventsourceflex183_trigger_filtered <= ((~irqarray11_interrupts[7]) & irqarray11_eventsourceflex183_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex183_trigger_filtered <= irqarray11_interrupts[7];
    end
end
assign irqarray11_eventsourceflex183_status = (irqarray11_interrupts[7] | irqarray11_trigger[7]);
always @(*) begin
    irqarray11_eventsourceflex184_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[8]) begin
        if (irqarray11_rising[8]) begin
            irqarray11_eventsourceflex184_trigger_filtered <= (irqarray11_interrupts[8] & (~irqarray11_eventsourceflex184_trigger_d));
        end else begin
            irqarray11_eventsourceflex184_trigger_filtered <= ((~irqarray11_interrupts[8]) & irqarray11_eventsourceflex184_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex184_trigger_filtered <= irqarray11_interrupts[8];
    end
end
assign irqarray11_eventsourceflex184_status = (irqarray11_interrupts[8] | irqarray11_trigger[8]);
always @(*) begin
    irqarray11_eventsourceflex185_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[9]) begin
        if (irqarray11_rising[9]) begin
            irqarray11_eventsourceflex185_trigger_filtered <= (irqarray11_interrupts[9] & (~irqarray11_eventsourceflex185_trigger_d));
        end else begin
            irqarray11_eventsourceflex185_trigger_filtered <= ((~irqarray11_interrupts[9]) & irqarray11_eventsourceflex185_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex185_trigger_filtered <= irqarray11_interrupts[9];
    end
end
assign irqarray11_eventsourceflex185_status = (irqarray11_interrupts[9] | irqarray11_trigger[9]);
always @(*) begin
    irqarray11_eventsourceflex186_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[10]) begin
        if (irqarray11_rising[10]) begin
            irqarray11_eventsourceflex186_trigger_filtered <= (irqarray11_interrupts[10] & (~irqarray11_eventsourceflex186_trigger_d));
        end else begin
            irqarray11_eventsourceflex186_trigger_filtered <= ((~irqarray11_interrupts[10]) & irqarray11_eventsourceflex186_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex186_trigger_filtered <= irqarray11_interrupts[10];
    end
end
assign irqarray11_eventsourceflex186_status = (irqarray11_interrupts[10] | irqarray11_trigger[10]);
always @(*) begin
    irqarray11_eventsourceflex187_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[11]) begin
        if (irqarray11_rising[11]) begin
            irqarray11_eventsourceflex187_trigger_filtered <= (irqarray11_interrupts[11] & (~irqarray11_eventsourceflex187_trigger_d));
        end else begin
            irqarray11_eventsourceflex187_trigger_filtered <= ((~irqarray11_interrupts[11]) & irqarray11_eventsourceflex187_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex187_trigger_filtered <= irqarray11_interrupts[11];
    end
end
assign irqarray11_eventsourceflex187_status = (irqarray11_interrupts[11] | irqarray11_trigger[11]);
always @(*) begin
    irqarray11_eventsourceflex188_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[12]) begin
        if (irqarray11_rising[12]) begin
            irqarray11_eventsourceflex188_trigger_filtered <= (irqarray11_interrupts[12] & (~irqarray11_eventsourceflex188_trigger_d));
        end else begin
            irqarray11_eventsourceflex188_trigger_filtered <= ((~irqarray11_interrupts[12]) & irqarray11_eventsourceflex188_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex188_trigger_filtered <= irqarray11_interrupts[12];
    end
end
assign irqarray11_eventsourceflex188_status = (irqarray11_interrupts[12] | irqarray11_trigger[12]);
always @(*) begin
    irqarray11_eventsourceflex189_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[13]) begin
        if (irqarray11_rising[13]) begin
            irqarray11_eventsourceflex189_trigger_filtered <= (irqarray11_interrupts[13] & (~irqarray11_eventsourceflex189_trigger_d));
        end else begin
            irqarray11_eventsourceflex189_trigger_filtered <= ((~irqarray11_interrupts[13]) & irqarray11_eventsourceflex189_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex189_trigger_filtered <= irqarray11_interrupts[13];
    end
end
assign irqarray11_eventsourceflex189_status = (irqarray11_interrupts[13] | irqarray11_trigger[13]);
always @(*) begin
    irqarray11_eventsourceflex190_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[14]) begin
        if (irqarray11_rising[14]) begin
            irqarray11_eventsourceflex190_trigger_filtered <= (irqarray11_interrupts[14] & (~irqarray11_eventsourceflex190_trigger_d));
        end else begin
            irqarray11_eventsourceflex190_trigger_filtered <= ((~irqarray11_interrupts[14]) & irqarray11_eventsourceflex190_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex190_trigger_filtered <= irqarray11_interrupts[14];
    end
end
assign irqarray11_eventsourceflex190_status = (irqarray11_interrupts[14] | irqarray11_trigger[14]);
always @(*) begin
    irqarray11_eventsourceflex191_trigger_filtered <= 1'd0;
    if (irqarray11_use_edge[15]) begin
        if (irqarray11_rising[15]) begin
            irqarray11_eventsourceflex191_trigger_filtered <= (irqarray11_interrupts[15] & (~irqarray11_eventsourceflex191_trigger_d));
        end else begin
            irqarray11_eventsourceflex191_trigger_filtered <= ((~irqarray11_interrupts[15]) & irqarray11_eventsourceflex191_trigger_d);
        end
    end else begin
        irqarray11_eventsourceflex191_trigger_filtered <= irqarray11_interrupts[15];
    end
end
assign irqarray11_eventsourceflex191_status = (irqarray11_interrupts[15] | irqarray11_trigger[15]);
assign irqarray12_interrupts = irq_remap12;
assign irqarray12_nc_b12s00 = irqarray12_eventsourceflex192_status;
assign irqarray12_nc_b12s01 = irqarray12_eventsourceflex192_pending;
always @(*) begin
    irqarray12_eventsourceflex192_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[0])) begin
        irqarray12_eventsourceflex192_clear <= 1'd1;
    end
end
assign irqarray12_nc_b12s10 = irqarray12_eventsourceflex193_status;
assign irqarray12_nc_b12s11 = irqarray12_eventsourceflex193_pending;
always @(*) begin
    irqarray12_eventsourceflex193_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[1])) begin
        irqarray12_eventsourceflex193_clear <= 1'd1;
    end
end
assign irqarray12_nc_b12s20 = irqarray12_eventsourceflex194_status;
assign irqarray12_nc_b12s21 = irqarray12_eventsourceflex194_pending;
always @(*) begin
    irqarray12_eventsourceflex194_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[2])) begin
        irqarray12_eventsourceflex194_clear <= 1'd1;
    end
end
assign irqarray12_nc_b12s30 = irqarray12_eventsourceflex195_status;
assign irqarray12_nc_b12s31 = irqarray12_eventsourceflex195_pending;
always @(*) begin
    irqarray12_eventsourceflex195_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[3])) begin
        irqarray12_eventsourceflex195_clear <= 1'd1;
    end
end
assign irqarray12_nc_b12s40 = irqarray12_eventsourceflex196_status;
assign irqarray12_nc_b12s41 = irqarray12_eventsourceflex196_pending;
always @(*) begin
    irqarray12_eventsourceflex196_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[4])) begin
        irqarray12_eventsourceflex196_clear <= 1'd1;
    end
end
assign irqarray12_nc_b12s50 = irqarray12_eventsourceflex197_status;
assign irqarray12_nc_b12s51 = irqarray12_eventsourceflex197_pending;
always @(*) begin
    irqarray12_eventsourceflex197_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[5])) begin
        irqarray12_eventsourceflex197_clear <= 1'd1;
    end
end
assign irqarray12_nc_b12s60 = irqarray12_eventsourceflex198_status;
assign irqarray12_nc_b12s61 = irqarray12_eventsourceflex198_pending;
always @(*) begin
    irqarray12_eventsourceflex198_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[6])) begin
        irqarray12_eventsourceflex198_clear <= 1'd1;
    end
end
assign irqarray12_nc_b12s70 = irqarray12_eventsourceflex199_status;
assign irqarray12_nc_b12s71 = irqarray12_eventsourceflex199_pending;
always @(*) begin
    irqarray12_eventsourceflex199_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[7])) begin
        irqarray12_eventsourceflex199_clear <= 1'd1;
    end
end
assign irqarray12_i2c0_nack0 = irqarray12_eventsourceflex200_status;
assign irqarray12_i2c0_nack1 = irqarray12_eventsourceflex200_pending;
always @(*) begin
    irqarray12_eventsourceflex200_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[8])) begin
        irqarray12_eventsourceflex200_clear <= 1'd1;
    end
end
assign irqarray12_i2c1_nack0 = irqarray12_eventsourceflex201_status;
assign irqarray12_i2c1_nack1 = irqarray12_eventsourceflex201_pending;
always @(*) begin
    irqarray12_eventsourceflex201_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[9])) begin
        irqarray12_eventsourceflex201_clear <= 1'd1;
    end
end
assign irqarray12_i2c2_nack0 = irqarray12_eventsourceflex202_status;
assign irqarray12_i2c2_nack1 = irqarray12_eventsourceflex202_pending;
always @(*) begin
    irqarray12_eventsourceflex202_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[10])) begin
        irqarray12_eventsourceflex202_clear <= 1'd1;
    end
end
assign irqarray12_i2c3_nack0 = irqarray12_eventsourceflex203_status;
assign irqarray12_i2c3_nack1 = irqarray12_eventsourceflex203_pending;
always @(*) begin
    irqarray12_eventsourceflex203_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[11])) begin
        irqarray12_eventsourceflex203_clear <= 1'd1;
    end
end
assign irqarray12_i2c0_err0 = irqarray12_eventsourceflex204_status;
assign irqarray12_i2c0_err1 = irqarray12_eventsourceflex204_pending;
always @(*) begin
    irqarray12_eventsourceflex204_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[12])) begin
        irqarray12_eventsourceflex204_clear <= 1'd1;
    end
end
assign irqarray12_i2c1_err0 = irqarray12_eventsourceflex205_status;
assign irqarray12_i2c1_err1 = irqarray12_eventsourceflex205_pending;
always @(*) begin
    irqarray12_eventsourceflex205_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[13])) begin
        irqarray12_eventsourceflex205_clear <= 1'd1;
    end
end
assign irqarray12_i2c2_err0 = irqarray12_eventsourceflex206_status;
assign irqarray12_i2c2_err1 = irqarray12_eventsourceflex206_pending;
always @(*) begin
    irqarray12_eventsourceflex206_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[14])) begin
        irqarray12_eventsourceflex206_clear <= 1'd1;
    end
end
assign irqarray12_i2c3_err0 = irqarray12_eventsourceflex207_status;
assign irqarray12_i2c3_err1 = irqarray12_eventsourceflex207_pending;
always @(*) begin
    irqarray12_eventsourceflex207_clear <= 1'd0;
    if ((irqarray12_pending_re & irqarray12_pending_r[15])) begin
        irqarray12_eventsourceflex207_clear <= 1'd1;
    end
end
assign irqarray12_irq = ((((((((((((((((irqarray12_pending_status[0] & irqarray12_enable_storage[0]) | (irqarray12_pending_status[1] & irqarray12_enable_storage[1])) | (irqarray12_pending_status[2] & irqarray12_enable_storage[2])) | (irqarray12_pending_status[3] & irqarray12_enable_storage[3])) | (irqarray12_pending_status[4] & irqarray12_enable_storage[4])) | (irqarray12_pending_status[5] & irqarray12_enable_storage[5])) | (irqarray12_pending_status[6] & irqarray12_enable_storage[6])) | (irqarray12_pending_status[7] & irqarray12_enable_storage[7])) | (irqarray12_pending_status[8] & irqarray12_enable_storage[8])) | (irqarray12_pending_status[9] & irqarray12_enable_storage[9])) | (irqarray12_pending_status[10] & irqarray12_enable_storage[10])) | (irqarray12_pending_status[11] & irqarray12_enable_storage[11])) | (irqarray12_pending_status[12] & irqarray12_enable_storage[12])) | (irqarray12_pending_status[13] & irqarray12_enable_storage[13])) | (irqarray12_pending_status[14] & irqarray12_enable_storage[14])) | (irqarray12_pending_status[15] & irqarray12_enable_storage[15]));
always @(*) begin
    irqarray12_eventsourceflex192_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[0]) begin
        if (irqarray12_rising[0]) begin
            irqarray12_eventsourceflex192_trigger_filtered <= (irqarray12_interrupts[0] & (~irqarray12_eventsourceflex192_trigger_d));
        end else begin
            irqarray12_eventsourceflex192_trigger_filtered <= ((~irqarray12_interrupts[0]) & irqarray12_eventsourceflex192_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex192_trigger_filtered <= irqarray12_interrupts[0];
    end
end
assign irqarray12_eventsourceflex192_status = (irqarray12_interrupts[0] | irqarray12_trigger[0]);
always @(*) begin
    irqarray12_eventsourceflex193_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[1]) begin
        if (irqarray12_rising[1]) begin
            irqarray12_eventsourceflex193_trigger_filtered <= (irqarray12_interrupts[1] & (~irqarray12_eventsourceflex193_trigger_d));
        end else begin
            irqarray12_eventsourceflex193_trigger_filtered <= ((~irqarray12_interrupts[1]) & irqarray12_eventsourceflex193_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex193_trigger_filtered <= irqarray12_interrupts[1];
    end
end
assign irqarray12_eventsourceflex193_status = (irqarray12_interrupts[1] | irqarray12_trigger[1]);
always @(*) begin
    irqarray12_eventsourceflex194_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[2]) begin
        if (irqarray12_rising[2]) begin
            irqarray12_eventsourceflex194_trigger_filtered <= (irqarray12_interrupts[2] & (~irqarray12_eventsourceflex194_trigger_d));
        end else begin
            irqarray12_eventsourceflex194_trigger_filtered <= ((~irqarray12_interrupts[2]) & irqarray12_eventsourceflex194_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex194_trigger_filtered <= irqarray12_interrupts[2];
    end
end
assign irqarray12_eventsourceflex194_status = (irqarray12_interrupts[2] | irqarray12_trigger[2]);
always @(*) begin
    irqarray12_eventsourceflex195_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[3]) begin
        if (irqarray12_rising[3]) begin
            irqarray12_eventsourceflex195_trigger_filtered <= (irqarray12_interrupts[3] & (~irqarray12_eventsourceflex195_trigger_d));
        end else begin
            irqarray12_eventsourceflex195_trigger_filtered <= ((~irqarray12_interrupts[3]) & irqarray12_eventsourceflex195_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex195_trigger_filtered <= irqarray12_interrupts[3];
    end
end
assign irqarray12_eventsourceflex195_status = (irqarray12_interrupts[3] | irqarray12_trigger[3]);
always @(*) begin
    irqarray12_eventsourceflex196_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[4]) begin
        if (irqarray12_rising[4]) begin
            irqarray12_eventsourceflex196_trigger_filtered <= (irqarray12_interrupts[4] & (~irqarray12_eventsourceflex196_trigger_d));
        end else begin
            irqarray12_eventsourceflex196_trigger_filtered <= ((~irqarray12_interrupts[4]) & irqarray12_eventsourceflex196_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex196_trigger_filtered <= irqarray12_interrupts[4];
    end
end
assign irqarray12_eventsourceflex196_status = (irqarray12_interrupts[4] | irqarray12_trigger[4]);
always @(*) begin
    irqarray12_eventsourceflex197_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[5]) begin
        if (irqarray12_rising[5]) begin
            irqarray12_eventsourceflex197_trigger_filtered <= (irqarray12_interrupts[5] & (~irqarray12_eventsourceflex197_trigger_d));
        end else begin
            irqarray12_eventsourceflex197_trigger_filtered <= ((~irqarray12_interrupts[5]) & irqarray12_eventsourceflex197_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex197_trigger_filtered <= irqarray12_interrupts[5];
    end
end
assign irqarray12_eventsourceflex197_status = (irqarray12_interrupts[5] | irqarray12_trigger[5]);
always @(*) begin
    irqarray12_eventsourceflex198_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[6]) begin
        if (irqarray12_rising[6]) begin
            irqarray12_eventsourceflex198_trigger_filtered <= (irqarray12_interrupts[6] & (~irqarray12_eventsourceflex198_trigger_d));
        end else begin
            irqarray12_eventsourceflex198_trigger_filtered <= ((~irqarray12_interrupts[6]) & irqarray12_eventsourceflex198_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex198_trigger_filtered <= irqarray12_interrupts[6];
    end
end
assign irqarray12_eventsourceflex198_status = (irqarray12_interrupts[6] | irqarray12_trigger[6]);
always @(*) begin
    irqarray12_eventsourceflex199_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[7]) begin
        if (irqarray12_rising[7]) begin
            irqarray12_eventsourceflex199_trigger_filtered <= (irqarray12_interrupts[7] & (~irqarray12_eventsourceflex199_trigger_d));
        end else begin
            irqarray12_eventsourceflex199_trigger_filtered <= ((~irqarray12_interrupts[7]) & irqarray12_eventsourceflex199_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex199_trigger_filtered <= irqarray12_interrupts[7];
    end
end
assign irqarray12_eventsourceflex199_status = (irqarray12_interrupts[7] | irqarray12_trigger[7]);
always @(*) begin
    irqarray12_eventsourceflex200_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[8]) begin
        if (irqarray12_rising[8]) begin
            irqarray12_eventsourceflex200_trigger_filtered <= (irqarray12_interrupts[8] & (~irqarray12_eventsourceflex200_trigger_d));
        end else begin
            irqarray12_eventsourceflex200_trigger_filtered <= ((~irqarray12_interrupts[8]) & irqarray12_eventsourceflex200_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex200_trigger_filtered <= irqarray12_interrupts[8];
    end
end
assign irqarray12_eventsourceflex200_status = (irqarray12_interrupts[8] | irqarray12_trigger[8]);
always @(*) begin
    irqarray12_eventsourceflex201_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[9]) begin
        if (irqarray12_rising[9]) begin
            irqarray12_eventsourceflex201_trigger_filtered <= (irqarray12_interrupts[9] & (~irqarray12_eventsourceflex201_trigger_d));
        end else begin
            irqarray12_eventsourceflex201_trigger_filtered <= ((~irqarray12_interrupts[9]) & irqarray12_eventsourceflex201_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex201_trigger_filtered <= irqarray12_interrupts[9];
    end
end
assign irqarray12_eventsourceflex201_status = (irqarray12_interrupts[9] | irqarray12_trigger[9]);
always @(*) begin
    irqarray12_eventsourceflex202_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[10]) begin
        if (irqarray12_rising[10]) begin
            irqarray12_eventsourceflex202_trigger_filtered <= (irqarray12_interrupts[10] & (~irqarray12_eventsourceflex202_trigger_d));
        end else begin
            irqarray12_eventsourceflex202_trigger_filtered <= ((~irqarray12_interrupts[10]) & irqarray12_eventsourceflex202_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex202_trigger_filtered <= irqarray12_interrupts[10];
    end
end
assign irqarray12_eventsourceflex202_status = (irqarray12_interrupts[10] | irqarray12_trigger[10]);
always @(*) begin
    irqarray12_eventsourceflex203_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[11]) begin
        if (irqarray12_rising[11]) begin
            irqarray12_eventsourceflex203_trigger_filtered <= (irqarray12_interrupts[11] & (~irqarray12_eventsourceflex203_trigger_d));
        end else begin
            irqarray12_eventsourceflex203_trigger_filtered <= ((~irqarray12_interrupts[11]) & irqarray12_eventsourceflex203_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex203_trigger_filtered <= irqarray12_interrupts[11];
    end
end
assign irqarray12_eventsourceflex203_status = (irqarray12_interrupts[11] | irqarray12_trigger[11]);
always @(*) begin
    irqarray12_eventsourceflex204_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[12]) begin
        if (irqarray12_rising[12]) begin
            irqarray12_eventsourceflex204_trigger_filtered <= (irqarray12_interrupts[12] & (~irqarray12_eventsourceflex204_trigger_d));
        end else begin
            irqarray12_eventsourceflex204_trigger_filtered <= ((~irqarray12_interrupts[12]) & irqarray12_eventsourceflex204_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex204_trigger_filtered <= irqarray12_interrupts[12];
    end
end
assign irqarray12_eventsourceflex204_status = (irqarray12_interrupts[12] | irqarray12_trigger[12]);
always @(*) begin
    irqarray12_eventsourceflex205_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[13]) begin
        if (irqarray12_rising[13]) begin
            irqarray12_eventsourceflex205_trigger_filtered <= (irqarray12_interrupts[13] & (~irqarray12_eventsourceflex205_trigger_d));
        end else begin
            irqarray12_eventsourceflex205_trigger_filtered <= ((~irqarray12_interrupts[13]) & irqarray12_eventsourceflex205_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex205_trigger_filtered <= irqarray12_interrupts[13];
    end
end
assign irqarray12_eventsourceflex205_status = (irqarray12_interrupts[13] | irqarray12_trigger[13]);
always @(*) begin
    irqarray12_eventsourceflex206_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[14]) begin
        if (irqarray12_rising[14]) begin
            irqarray12_eventsourceflex206_trigger_filtered <= (irqarray12_interrupts[14] & (~irqarray12_eventsourceflex206_trigger_d));
        end else begin
            irqarray12_eventsourceflex206_trigger_filtered <= ((~irqarray12_interrupts[14]) & irqarray12_eventsourceflex206_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex206_trigger_filtered <= irqarray12_interrupts[14];
    end
end
assign irqarray12_eventsourceflex206_status = (irqarray12_interrupts[14] | irqarray12_trigger[14]);
always @(*) begin
    irqarray12_eventsourceflex207_trigger_filtered <= 1'd0;
    if (irqarray12_use_edge[15]) begin
        if (irqarray12_rising[15]) begin
            irqarray12_eventsourceflex207_trigger_filtered <= (irqarray12_interrupts[15] & (~irqarray12_eventsourceflex207_trigger_d));
        end else begin
            irqarray12_eventsourceflex207_trigger_filtered <= ((~irqarray12_interrupts[15]) & irqarray12_eventsourceflex207_trigger_d);
        end
    end else begin
        irqarray12_eventsourceflex207_trigger_filtered <= irqarray12_interrupts[15];
    end
end
assign irqarray12_eventsourceflex207_status = (irqarray12_interrupts[15] | irqarray12_trigger[15]);
assign irqarray13_interrupts = irq_remap13;
assign irqarray13_coresuberr0 = irqarray13_eventsourceflex208_status;
assign irqarray13_coresuberr1 = irqarray13_eventsourceflex208_pending;
always @(*) begin
    irqarray13_eventsourceflex208_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[0])) begin
        irqarray13_eventsourceflex208_clear <= 1'd1;
    end
end
assign irqarray13_sceerr0 = irqarray13_eventsourceflex209_status;
assign irqarray13_sceerr1 = irqarray13_eventsourceflex209_pending;
always @(*) begin
    irqarray13_eventsourceflex209_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[1])) begin
        irqarray13_eventsourceflex209_clear <= 1'd1;
    end
end
assign irqarray13_ifsuberr0 = irqarray13_eventsourceflex210_status;
assign irqarray13_ifsuberr1 = irqarray13_eventsourceflex210_pending;
always @(*) begin
    irqarray13_eventsourceflex210_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[2])) begin
        irqarray13_eventsourceflex210_clear <= 1'd1;
    end
end
assign irqarray13_secirq0 = irqarray13_eventsourceflex211_status;
assign irqarray13_secirq1 = irqarray13_eventsourceflex211_pending;
always @(*) begin
    irqarray13_eventsourceflex211_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[3])) begin
        irqarray13_eventsourceflex211_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s40 = irqarray13_eventsourceflex212_status;
assign irqarray13_nc_b13s41 = irqarray13_eventsourceflex212_pending;
always @(*) begin
    irqarray13_eventsourceflex212_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[4])) begin
        irqarray13_eventsourceflex212_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s50 = irqarray13_eventsourceflex213_status;
assign irqarray13_nc_b13s51 = irqarray13_eventsourceflex213_pending;
always @(*) begin
    irqarray13_eventsourceflex213_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[5])) begin
        irqarray13_eventsourceflex213_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s60 = irqarray13_eventsourceflex214_status;
assign irqarray13_nc_b13s61 = irqarray13_eventsourceflex214_pending;
always @(*) begin
    irqarray13_eventsourceflex214_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[6])) begin
        irqarray13_eventsourceflex214_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s70 = irqarray13_eventsourceflex215_status;
assign irqarray13_nc_b13s71 = irqarray13_eventsourceflex215_pending;
always @(*) begin
    irqarray13_eventsourceflex215_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[7])) begin
        irqarray13_eventsourceflex215_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s80 = irqarray13_eventsourceflex216_status;
assign irqarray13_nc_b13s81 = irqarray13_eventsourceflex216_pending;
always @(*) begin
    irqarray13_eventsourceflex216_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[8])) begin
        irqarray13_eventsourceflex216_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s90 = irqarray13_eventsourceflex217_status;
assign irqarray13_nc_b13s91 = irqarray13_eventsourceflex217_pending;
always @(*) begin
    irqarray13_eventsourceflex217_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[9])) begin
        irqarray13_eventsourceflex217_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s100 = irqarray13_eventsourceflex218_status;
assign irqarray13_nc_b13s101 = irqarray13_eventsourceflex218_pending;
always @(*) begin
    irqarray13_eventsourceflex218_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[10])) begin
        irqarray13_eventsourceflex218_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s110 = irqarray13_eventsourceflex219_status;
assign irqarray13_nc_b13s111 = irqarray13_eventsourceflex219_pending;
always @(*) begin
    irqarray13_eventsourceflex219_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[11])) begin
        irqarray13_eventsourceflex219_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s120 = irqarray13_eventsourceflex220_status;
assign irqarray13_nc_b13s121 = irqarray13_eventsourceflex220_pending;
always @(*) begin
    irqarray13_eventsourceflex220_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[12])) begin
        irqarray13_eventsourceflex220_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s130 = irqarray13_eventsourceflex221_status;
assign irqarray13_nc_b13s131 = irqarray13_eventsourceflex221_pending;
always @(*) begin
    irqarray13_eventsourceflex221_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[13])) begin
        irqarray13_eventsourceflex221_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s140 = irqarray13_eventsourceflex222_status;
assign irqarray13_nc_b13s141 = irqarray13_eventsourceflex222_pending;
always @(*) begin
    irqarray13_eventsourceflex222_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[14])) begin
        irqarray13_eventsourceflex222_clear <= 1'd1;
    end
end
assign irqarray13_nc_b13s150 = irqarray13_eventsourceflex223_status;
assign irqarray13_nc_b13s151 = irqarray13_eventsourceflex223_pending;
always @(*) begin
    irqarray13_eventsourceflex223_clear <= 1'd0;
    if ((irqarray13_pending_re & irqarray13_pending_r[15])) begin
        irqarray13_eventsourceflex223_clear <= 1'd1;
    end
end
assign irqarray13_irq = ((((((((((((((((irqarray13_pending_status[0] & irqarray13_enable_storage[0]) | (irqarray13_pending_status[1] & irqarray13_enable_storage[1])) | (irqarray13_pending_status[2] & irqarray13_enable_storage[2])) | (irqarray13_pending_status[3] & irqarray13_enable_storage[3])) | (irqarray13_pending_status[4] & irqarray13_enable_storage[4])) | (irqarray13_pending_status[5] & irqarray13_enable_storage[5])) | (irqarray13_pending_status[6] & irqarray13_enable_storage[6])) | (irqarray13_pending_status[7] & irqarray13_enable_storage[7])) | (irqarray13_pending_status[8] & irqarray13_enable_storage[8])) | (irqarray13_pending_status[9] & irqarray13_enable_storage[9])) | (irqarray13_pending_status[10] & irqarray13_enable_storage[10])) | (irqarray13_pending_status[11] & irqarray13_enable_storage[11])) | (irqarray13_pending_status[12] & irqarray13_enable_storage[12])) | (irqarray13_pending_status[13] & irqarray13_enable_storage[13])) | (irqarray13_pending_status[14] & irqarray13_enable_storage[14])) | (irqarray13_pending_status[15] & irqarray13_enable_storage[15]));
always @(*) begin
    irqarray13_eventsourceflex208_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[0]) begin
        if (irqarray13_rising[0]) begin
            irqarray13_eventsourceflex208_trigger_filtered <= (irqarray13_interrupts[0] & (~irqarray13_eventsourceflex208_trigger_d));
        end else begin
            irqarray13_eventsourceflex208_trigger_filtered <= ((~irqarray13_interrupts[0]) & irqarray13_eventsourceflex208_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex208_trigger_filtered <= irqarray13_interrupts[0];
    end
end
assign irqarray13_eventsourceflex208_status = (irqarray13_interrupts[0] | irqarray13_trigger[0]);
always @(*) begin
    irqarray13_eventsourceflex209_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[1]) begin
        if (irqarray13_rising[1]) begin
            irqarray13_eventsourceflex209_trigger_filtered <= (irqarray13_interrupts[1] & (~irqarray13_eventsourceflex209_trigger_d));
        end else begin
            irqarray13_eventsourceflex209_trigger_filtered <= ((~irqarray13_interrupts[1]) & irqarray13_eventsourceflex209_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex209_trigger_filtered <= irqarray13_interrupts[1];
    end
end
assign irqarray13_eventsourceflex209_status = (irqarray13_interrupts[1] | irqarray13_trigger[1]);
always @(*) begin
    irqarray13_eventsourceflex210_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[2]) begin
        if (irqarray13_rising[2]) begin
            irqarray13_eventsourceflex210_trigger_filtered <= (irqarray13_interrupts[2] & (~irqarray13_eventsourceflex210_trigger_d));
        end else begin
            irqarray13_eventsourceflex210_trigger_filtered <= ((~irqarray13_interrupts[2]) & irqarray13_eventsourceflex210_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex210_trigger_filtered <= irqarray13_interrupts[2];
    end
end
assign irqarray13_eventsourceflex210_status = (irqarray13_interrupts[2] | irqarray13_trigger[2]);
always @(*) begin
    irqarray13_eventsourceflex211_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[3]) begin
        if (irqarray13_rising[3]) begin
            irqarray13_eventsourceflex211_trigger_filtered <= (irqarray13_interrupts[3] & (~irqarray13_eventsourceflex211_trigger_d));
        end else begin
            irqarray13_eventsourceflex211_trigger_filtered <= ((~irqarray13_interrupts[3]) & irqarray13_eventsourceflex211_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex211_trigger_filtered <= irqarray13_interrupts[3];
    end
end
assign irqarray13_eventsourceflex211_status = (irqarray13_interrupts[3] | irqarray13_trigger[3]);
always @(*) begin
    irqarray13_eventsourceflex212_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[4]) begin
        if (irqarray13_rising[4]) begin
            irqarray13_eventsourceflex212_trigger_filtered <= (irqarray13_interrupts[4] & (~irqarray13_eventsourceflex212_trigger_d));
        end else begin
            irqarray13_eventsourceflex212_trigger_filtered <= ((~irqarray13_interrupts[4]) & irqarray13_eventsourceflex212_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex212_trigger_filtered <= irqarray13_interrupts[4];
    end
end
assign irqarray13_eventsourceflex212_status = (irqarray13_interrupts[4] | irqarray13_trigger[4]);
always @(*) begin
    irqarray13_eventsourceflex213_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[5]) begin
        if (irqarray13_rising[5]) begin
            irqarray13_eventsourceflex213_trigger_filtered <= (irqarray13_interrupts[5] & (~irqarray13_eventsourceflex213_trigger_d));
        end else begin
            irqarray13_eventsourceflex213_trigger_filtered <= ((~irqarray13_interrupts[5]) & irqarray13_eventsourceflex213_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex213_trigger_filtered <= irqarray13_interrupts[5];
    end
end
assign irqarray13_eventsourceflex213_status = (irqarray13_interrupts[5] | irqarray13_trigger[5]);
always @(*) begin
    irqarray13_eventsourceflex214_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[6]) begin
        if (irqarray13_rising[6]) begin
            irqarray13_eventsourceflex214_trigger_filtered <= (irqarray13_interrupts[6] & (~irqarray13_eventsourceflex214_trigger_d));
        end else begin
            irqarray13_eventsourceflex214_trigger_filtered <= ((~irqarray13_interrupts[6]) & irqarray13_eventsourceflex214_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex214_trigger_filtered <= irqarray13_interrupts[6];
    end
end
assign irqarray13_eventsourceflex214_status = (irqarray13_interrupts[6] | irqarray13_trigger[6]);
always @(*) begin
    irqarray13_eventsourceflex215_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[7]) begin
        if (irqarray13_rising[7]) begin
            irqarray13_eventsourceflex215_trigger_filtered <= (irqarray13_interrupts[7] & (~irqarray13_eventsourceflex215_trigger_d));
        end else begin
            irqarray13_eventsourceflex215_trigger_filtered <= ((~irqarray13_interrupts[7]) & irqarray13_eventsourceflex215_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex215_trigger_filtered <= irqarray13_interrupts[7];
    end
end
assign irqarray13_eventsourceflex215_status = (irqarray13_interrupts[7] | irqarray13_trigger[7]);
always @(*) begin
    irqarray13_eventsourceflex216_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[8]) begin
        if (irqarray13_rising[8]) begin
            irqarray13_eventsourceflex216_trigger_filtered <= (irqarray13_interrupts[8] & (~irqarray13_eventsourceflex216_trigger_d));
        end else begin
            irqarray13_eventsourceflex216_trigger_filtered <= ((~irqarray13_interrupts[8]) & irqarray13_eventsourceflex216_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex216_trigger_filtered <= irqarray13_interrupts[8];
    end
end
assign irqarray13_eventsourceflex216_status = (irqarray13_interrupts[8] | irqarray13_trigger[8]);
always @(*) begin
    irqarray13_eventsourceflex217_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[9]) begin
        if (irqarray13_rising[9]) begin
            irqarray13_eventsourceflex217_trigger_filtered <= (irqarray13_interrupts[9] & (~irqarray13_eventsourceflex217_trigger_d));
        end else begin
            irqarray13_eventsourceflex217_trigger_filtered <= ((~irqarray13_interrupts[9]) & irqarray13_eventsourceflex217_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex217_trigger_filtered <= irqarray13_interrupts[9];
    end
end
assign irqarray13_eventsourceflex217_status = (irqarray13_interrupts[9] | irqarray13_trigger[9]);
always @(*) begin
    irqarray13_eventsourceflex218_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[10]) begin
        if (irqarray13_rising[10]) begin
            irqarray13_eventsourceflex218_trigger_filtered <= (irqarray13_interrupts[10] & (~irqarray13_eventsourceflex218_trigger_d));
        end else begin
            irqarray13_eventsourceflex218_trigger_filtered <= ((~irqarray13_interrupts[10]) & irqarray13_eventsourceflex218_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex218_trigger_filtered <= irqarray13_interrupts[10];
    end
end
assign irqarray13_eventsourceflex218_status = (irqarray13_interrupts[10] | irqarray13_trigger[10]);
always @(*) begin
    irqarray13_eventsourceflex219_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[11]) begin
        if (irqarray13_rising[11]) begin
            irqarray13_eventsourceflex219_trigger_filtered <= (irqarray13_interrupts[11] & (~irqarray13_eventsourceflex219_trigger_d));
        end else begin
            irqarray13_eventsourceflex219_trigger_filtered <= ((~irqarray13_interrupts[11]) & irqarray13_eventsourceflex219_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex219_trigger_filtered <= irqarray13_interrupts[11];
    end
end
assign irqarray13_eventsourceflex219_status = (irqarray13_interrupts[11] | irqarray13_trigger[11]);
always @(*) begin
    irqarray13_eventsourceflex220_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[12]) begin
        if (irqarray13_rising[12]) begin
            irqarray13_eventsourceflex220_trigger_filtered <= (irqarray13_interrupts[12] & (~irqarray13_eventsourceflex220_trigger_d));
        end else begin
            irqarray13_eventsourceflex220_trigger_filtered <= ((~irqarray13_interrupts[12]) & irqarray13_eventsourceflex220_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex220_trigger_filtered <= irqarray13_interrupts[12];
    end
end
assign irqarray13_eventsourceflex220_status = (irqarray13_interrupts[12] | irqarray13_trigger[12]);
always @(*) begin
    irqarray13_eventsourceflex221_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[13]) begin
        if (irqarray13_rising[13]) begin
            irqarray13_eventsourceflex221_trigger_filtered <= (irqarray13_interrupts[13] & (~irqarray13_eventsourceflex221_trigger_d));
        end else begin
            irqarray13_eventsourceflex221_trigger_filtered <= ((~irqarray13_interrupts[13]) & irqarray13_eventsourceflex221_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex221_trigger_filtered <= irqarray13_interrupts[13];
    end
end
assign irqarray13_eventsourceflex221_status = (irqarray13_interrupts[13] | irqarray13_trigger[13]);
always @(*) begin
    irqarray13_eventsourceflex222_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[14]) begin
        if (irqarray13_rising[14]) begin
            irqarray13_eventsourceflex222_trigger_filtered <= (irqarray13_interrupts[14] & (~irqarray13_eventsourceflex222_trigger_d));
        end else begin
            irqarray13_eventsourceflex222_trigger_filtered <= ((~irqarray13_interrupts[14]) & irqarray13_eventsourceflex222_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex222_trigger_filtered <= irqarray13_interrupts[14];
    end
end
assign irqarray13_eventsourceflex222_status = (irqarray13_interrupts[14] | irqarray13_trigger[14]);
always @(*) begin
    irqarray13_eventsourceflex223_trigger_filtered <= 1'd0;
    if (irqarray13_use_edge[15]) begin
        if (irqarray13_rising[15]) begin
            irqarray13_eventsourceflex223_trigger_filtered <= (irqarray13_interrupts[15] & (~irqarray13_eventsourceflex223_trigger_d));
        end else begin
            irqarray13_eventsourceflex223_trigger_filtered <= ((~irqarray13_interrupts[15]) & irqarray13_eventsourceflex223_trigger_d);
        end
    end else begin
        irqarray13_eventsourceflex223_trigger_filtered <= irqarray13_interrupts[15];
    end
end
assign irqarray13_eventsourceflex223_status = (irqarray13_interrupts[15] | irqarray13_trigger[15]);
assign irqarray14_interrupts = irq_remap14;
assign irqarray14_uart2_rx_dupe0 = irqarray14_eventsourceflex224_status;
assign irqarray14_uart2_rx_dupe1 = irqarray14_eventsourceflex224_pending;
always @(*) begin
    irqarray14_eventsourceflex224_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[0])) begin
        irqarray14_eventsourceflex224_clear <= 1'd1;
    end
end
assign irqarray14_uart2_tx_dupe0 = irqarray14_eventsourceflex225_status;
assign irqarray14_uart2_tx_dupe1 = irqarray14_eventsourceflex225_pending;
always @(*) begin
    irqarray14_eventsourceflex225_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[1])) begin
        irqarray14_eventsourceflex225_clear <= 1'd1;
    end
end
assign irqarray14_uart2_rx_char_dupe0 = irqarray14_eventsourceflex226_status;
assign irqarray14_uart2_rx_char_dupe1 = irqarray14_eventsourceflex226_pending;
always @(*) begin
    irqarray14_eventsourceflex226_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[2])) begin
        irqarray14_eventsourceflex226_clear <= 1'd1;
    end
end
assign irqarray14_uart2_err_dupe0 = irqarray14_eventsourceflex227_status;
assign irqarray14_uart2_err_dupe1 = irqarray14_eventsourceflex227_pending;
always @(*) begin
    irqarray14_eventsourceflex227_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[3])) begin
        irqarray14_eventsourceflex227_clear <= 1'd1;
    end
end
assign irqarray14_uart3_rx_dupe0 = irqarray14_eventsourceflex228_status;
assign irqarray14_uart3_rx_dupe1 = irqarray14_eventsourceflex228_pending;
always @(*) begin
    irqarray14_eventsourceflex228_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[4])) begin
        irqarray14_eventsourceflex228_clear <= 1'd1;
    end
end
assign irqarray14_uart3_tx_dupe0 = irqarray14_eventsourceflex229_status;
assign irqarray14_uart3_tx_dupe1 = irqarray14_eventsourceflex229_pending;
always @(*) begin
    irqarray14_eventsourceflex229_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[5])) begin
        irqarray14_eventsourceflex229_clear <= 1'd1;
    end
end
assign irqarray14_uart3_rx_char_dupe0 = irqarray14_eventsourceflex230_status;
assign irqarray14_uart3_rx_char_dupe1 = irqarray14_eventsourceflex230_pending;
always @(*) begin
    irqarray14_eventsourceflex230_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[6])) begin
        irqarray14_eventsourceflex230_clear <= 1'd1;
    end
end
assign irqarray14_uart3_err_dupe0 = irqarray14_eventsourceflex231_status;
assign irqarray14_uart3_err_dupe1 = irqarray14_eventsourceflex231_pending;
always @(*) begin
    irqarray14_eventsourceflex231_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[7])) begin
        irqarray14_eventsourceflex231_clear <= 1'd1;
    end
end
assign irqarray14_trng_done_dupe0 = irqarray14_eventsourceflex232_status;
assign irqarray14_trng_done_dupe1 = irqarray14_eventsourceflex232_pending;
always @(*) begin
    irqarray14_eventsourceflex232_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[8])) begin
        irqarray14_eventsourceflex232_clear <= 1'd1;
    end
end
assign irqarray14_nc_b14s90 = irqarray14_eventsourceflex233_status;
assign irqarray14_nc_b14s91 = irqarray14_eventsourceflex233_pending;
always @(*) begin
    irqarray14_eventsourceflex233_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[9])) begin
        irqarray14_eventsourceflex233_clear <= 1'd1;
    end
end
assign irqarray14_nc_b14s100 = irqarray14_eventsourceflex234_status;
assign irqarray14_nc_b14s101 = irqarray14_eventsourceflex234_pending;
always @(*) begin
    irqarray14_eventsourceflex234_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[10])) begin
        irqarray14_eventsourceflex234_clear <= 1'd1;
    end
end
assign irqarray14_nc_b14s110 = irqarray14_eventsourceflex235_status;
assign irqarray14_nc_b14s111 = irqarray14_eventsourceflex235_pending;
always @(*) begin
    irqarray14_eventsourceflex235_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[11])) begin
        irqarray14_eventsourceflex235_clear <= 1'd1;
    end
end
assign irqarray14_nc_b14s120 = irqarray14_eventsourceflex236_status;
assign irqarray14_nc_b14s121 = irqarray14_eventsourceflex236_pending;
always @(*) begin
    irqarray14_eventsourceflex236_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[12])) begin
        irqarray14_eventsourceflex236_clear <= 1'd1;
    end
end
assign irqarray14_nc_b14s130 = irqarray14_eventsourceflex237_status;
assign irqarray14_nc_b14s131 = irqarray14_eventsourceflex237_pending;
always @(*) begin
    irqarray14_eventsourceflex237_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[13])) begin
        irqarray14_eventsourceflex237_clear <= 1'd1;
    end
end
assign irqarray14_nc_b14s140 = irqarray14_eventsourceflex238_status;
assign irqarray14_nc_b14s141 = irqarray14_eventsourceflex238_pending;
always @(*) begin
    irqarray14_eventsourceflex238_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[14])) begin
        irqarray14_eventsourceflex238_clear <= 1'd1;
    end
end
assign irqarray14_nc_b14s150 = irqarray14_eventsourceflex239_status;
assign irqarray14_nc_b14s151 = irqarray14_eventsourceflex239_pending;
always @(*) begin
    irqarray14_eventsourceflex239_clear <= 1'd0;
    if ((irqarray14_pending_re & irqarray14_pending_r[15])) begin
        irqarray14_eventsourceflex239_clear <= 1'd1;
    end
end
assign irqarray14_irq = ((((((((((((((((irqarray14_pending_status[0] & irqarray14_enable_storage[0]) | (irqarray14_pending_status[1] & irqarray14_enable_storage[1])) | (irqarray14_pending_status[2] & irqarray14_enable_storage[2])) | (irqarray14_pending_status[3] & irqarray14_enable_storage[3])) | (irqarray14_pending_status[4] & irqarray14_enable_storage[4])) | (irqarray14_pending_status[5] & irqarray14_enable_storage[5])) | (irqarray14_pending_status[6] & irqarray14_enable_storage[6])) | (irqarray14_pending_status[7] & irqarray14_enable_storage[7])) | (irqarray14_pending_status[8] & irqarray14_enable_storage[8])) | (irqarray14_pending_status[9] & irqarray14_enable_storage[9])) | (irqarray14_pending_status[10] & irqarray14_enable_storage[10])) | (irqarray14_pending_status[11] & irqarray14_enable_storage[11])) | (irqarray14_pending_status[12] & irqarray14_enable_storage[12])) | (irqarray14_pending_status[13] & irqarray14_enable_storage[13])) | (irqarray14_pending_status[14] & irqarray14_enable_storage[14])) | (irqarray14_pending_status[15] & irqarray14_enable_storage[15]));
always @(*) begin
    irqarray14_eventsourceflex224_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[0]) begin
        if (irqarray14_rising[0]) begin
            irqarray14_eventsourceflex224_trigger_filtered <= (irqarray14_interrupts[0] & (~irqarray14_eventsourceflex224_trigger_d));
        end else begin
            irqarray14_eventsourceflex224_trigger_filtered <= ((~irqarray14_interrupts[0]) & irqarray14_eventsourceflex224_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex224_trigger_filtered <= irqarray14_interrupts[0];
    end
end
assign irqarray14_eventsourceflex224_status = (irqarray14_interrupts[0] | irqarray14_trigger[0]);
always @(*) begin
    irqarray14_eventsourceflex225_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[1]) begin
        if (irqarray14_rising[1]) begin
            irqarray14_eventsourceflex225_trigger_filtered <= (irqarray14_interrupts[1] & (~irqarray14_eventsourceflex225_trigger_d));
        end else begin
            irqarray14_eventsourceflex225_trigger_filtered <= ((~irqarray14_interrupts[1]) & irqarray14_eventsourceflex225_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex225_trigger_filtered <= irqarray14_interrupts[1];
    end
end
assign irqarray14_eventsourceflex225_status = (irqarray14_interrupts[1] | irqarray14_trigger[1]);
always @(*) begin
    irqarray14_eventsourceflex226_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[2]) begin
        if (irqarray14_rising[2]) begin
            irqarray14_eventsourceflex226_trigger_filtered <= (irqarray14_interrupts[2] & (~irqarray14_eventsourceflex226_trigger_d));
        end else begin
            irqarray14_eventsourceflex226_trigger_filtered <= ((~irqarray14_interrupts[2]) & irqarray14_eventsourceflex226_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex226_trigger_filtered <= irqarray14_interrupts[2];
    end
end
assign irqarray14_eventsourceflex226_status = (irqarray14_interrupts[2] | irqarray14_trigger[2]);
always @(*) begin
    irqarray14_eventsourceflex227_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[3]) begin
        if (irqarray14_rising[3]) begin
            irqarray14_eventsourceflex227_trigger_filtered <= (irqarray14_interrupts[3] & (~irqarray14_eventsourceflex227_trigger_d));
        end else begin
            irqarray14_eventsourceflex227_trigger_filtered <= ((~irqarray14_interrupts[3]) & irqarray14_eventsourceflex227_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex227_trigger_filtered <= irqarray14_interrupts[3];
    end
end
assign irqarray14_eventsourceflex227_status = (irqarray14_interrupts[3] | irqarray14_trigger[3]);
always @(*) begin
    irqarray14_eventsourceflex228_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[4]) begin
        if (irqarray14_rising[4]) begin
            irqarray14_eventsourceflex228_trigger_filtered <= (irqarray14_interrupts[4] & (~irqarray14_eventsourceflex228_trigger_d));
        end else begin
            irqarray14_eventsourceflex228_trigger_filtered <= ((~irqarray14_interrupts[4]) & irqarray14_eventsourceflex228_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex228_trigger_filtered <= irqarray14_interrupts[4];
    end
end
assign irqarray14_eventsourceflex228_status = (irqarray14_interrupts[4] | irqarray14_trigger[4]);
always @(*) begin
    irqarray14_eventsourceflex229_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[5]) begin
        if (irqarray14_rising[5]) begin
            irqarray14_eventsourceflex229_trigger_filtered <= (irqarray14_interrupts[5] & (~irqarray14_eventsourceflex229_trigger_d));
        end else begin
            irqarray14_eventsourceflex229_trigger_filtered <= ((~irqarray14_interrupts[5]) & irqarray14_eventsourceflex229_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex229_trigger_filtered <= irqarray14_interrupts[5];
    end
end
assign irqarray14_eventsourceflex229_status = (irqarray14_interrupts[5] | irqarray14_trigger[5]);
always @(*) begin
    irqarray14_eventsourceflex230_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[6]) begin
        if (irqarray14_rising[6]) begin
            irqarray14_eventsourceflex230_trigger_filtered <= (irqarray14_interrupts[6] & (~irqarray14_eventsourceflex230_trigger_d));
        end else begin
            irqarray14_eventsourceflex230_trigger_filtered <= ((~irqarray14_interrupts[6]) & irqarray14_eventsourceflex230_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex230_trigger_filtered <= irqarray14_interrupts[6];
    end
end
assign irqarray14_eventsourceflex230_status = (irqarray14_interrupts[6] | irqarray14_trigger[6]);
always @(*) begin
    irqarray14_eventsourceflex231_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[7]) begin
        if (irqarray14_rising[7]) begin
            irqarray14_eventsourceflex231_trigger_filtered <= (irqarray14_interrupts[7] & (~irqarray14_eventsourceflex231_trigger_d));
        end else begin
            irqarray14_eventsourceflex231_trigger_filtered <= ((~irqarray14_interrupts[7]) & irqarray14_eventsourceflex231_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex231_trigger_filtered <= irqarray14_interrupts[7];
    end
end
assign irqarray14_eventsourceflex231_status = (irqarray14_interrupts[7] | irqarray14_trigger[7]);
always @(*) begin
    irqarray14_eventsourceflex232_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[8]) begin
        if (irqarray14_rising[8]) begin
            irqarray14_eventsourceflex232_trigger_filtered <= (irqarray14_interrupts[8] & (~irqarray14_eventsourceflex232_trigger_d));
        end else begin
            irqarray14_eventsourceflex232_trigger_filtered <= ((~irqarray14_interrupts[8]) & irqarray14_eventsourceflex232_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex232_trigger_filtered <= irqarray14_interrupts[8];
    end
end
assign irqarray14_eventsourceflex232_status = (irqarray14_interrupts[8] | irqarray14_trigger[8]);
always @(*) begin
    irqarray14_eventsourceflex233_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[9]) begin
        if (irqarray14_rising[9]) begin
            irqarray14_eventsourceflex233_trigger_filtered <= (irqarray14_interrupts[9] & (~irqarray14_eventsourceflex233_trigger_d));
        end else begin
            irqarray14_eventsourceflex233_trigger_filtered <= ((~irqarray14_interrupts[9]) & irqarray14_eventsourceflex233_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex233_trigger_filtered <= irqarray14_interrupts[9];
    end
end
assign irqarray14_eventsourceflex233_status = (irqarray14_interrupts[9] | irqarray14_trigger[9]);
always @(*) begin
    irqarray14_eventsourceflex234_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[10]) begin
        if (irqarray14_rising[10]) begin
            irqarray14_eventsourceflex234_trigger_filtered <= (irqarray14_interrupts[10] & (~irqarray14_eventsourceflex234_trigger_d));
        end else begin
            irqarray14_eventsourceflex234_trigger_filtered <= ((~irqarray14_interrupts[10]) & irqarray14_eventsourceflex234_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex234_trigger_filtered <= irqarray14_interrupts[10];
    end
end
assign irqarray14_eventsourceflex234_status = (irqarray14_interrupts[10] | irqarray14_trigger[10]);
always @(*) begin
    irqarray14_eventsourceflex235_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[11]) begin
        if (irqarray14_rising[11]) begin
            irqarray14_eventsourceflex235_trigger_filtered <= (irqarray14_interrupts[11] & (~irqarray14_eventsourceflex235_trigger_d));
        end else begin
            irqarray14_eventsourceflex235_trigger_filtered <= ((~irqarray14_interrupts[11]) & irqarray14_eventsourceflex235_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex235_trigger_filtered <= irqarray14_interrupts[11];
    end
end
assign irqarray14_eventsourceflex235_status = (irqarray14_interrupts[11] | irqarray14_trigger[11]);
always @(*) begin
    irqarray14_eventsourceflex236_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[12]) begin
        if (irqarray14_rising[12]) begin
            irqarray14_eventsourceflex236_trigger_filtered <= (irqarray14_interrupts[12] & (~irqarray14_eventsourceflex236_trigger_d));
        end else begin
            irqarray14_eventsourceflex236_trigger_filtered <= ((~irqarray14_interrupts[12]) & irqarray14_eventsourceflex236_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex236_trigger_filtered <= irqarray14_interrupts[12];
    end
end
assign irqarray14_eventsourceflex236_status = (irqarray14_interrupts[12] | irqarray14_trigger[12]);
always @(*) begin
    irqarray14_eventsourceflex237_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[13]) begin
        if (irqarray14_rising[13]) begin
            irqarray14_eventsourceflex237_trigger_filtered <= (irqarray14_interrupts[13] & (~irqarray14_eventsourceflex237_trigger_d));
        end else begin
            irqarray14_eventsourceflex237_trigger_filtered <= ((~irqarray14_interrupts[13]) & irqarray14_eventsourceflex237_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex237_trigger_filtered <= irqarray14_interrupts[13];
    end
end
assign irqarray14_eventsourceflex237_status = (irqarray14_interrupts[13] | irqarray14_trigger[13]);
always @(*) begin
    irqarray14_eventsourceflex238_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[14]) begin
        if (irqarray14_rising[14]) begin
            irqarray14_eventsourceflex238_trigger_filtered <= (irqarray14_interrupts[14] & (~irqarray14_eventsourceflex238_trigger_d));
        end else begin
            irqarray14_eventsourceflex238_trigger_filtered <= ((~irqarray14_interrupts[14]) & irqarray14_eventsourceflex238_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex238_trigger_filtered <= irqarray14_interrupts[14];
    end
end
assign irqarray14_eventsourceflex238_status = (irqarray14_interrupts[14] | irqarray14_trigger[14]);
always @(*) begin
    irqarray14_eventsourceflex239_trigger_filtered <= 1'd0;
    if (irqarray14_use_edge[15]) begin
        if (irqarray14_rising[15]) begin
            irqarray14_eventsourceflex239_trigger_filtered <= (irqarray14_interrupts[15] & (~irqarray14_eventsourceflex239_trigger_d));
        end else begin
            irqarray14_eventsourceflex239_trigger_filtered <= ((~irqarray14_interrupts[15]) & irqarray14_eventsourceflex239_trigger_d);
        end
    end else begin
        irqarray14_eventsourceflex239_trigger_filtered <= irqarray14_interrupts[15];
    end
end
assign irqarray14_eventsourceflex239_status = (irqarray14_interrupts[15] | irqarray14_trigger[15]);
assign irqarray15_interrupts = irq_remap15;
assign irqarray15_sec00 = irqarray15_eventsourceflex240_status;
assign irqarray15_sec01 = irqarray15_eventsourceflex240_pending;
always @(*) begin
    irqarray15_eventsourceflex240_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[0])) begin
        irqarray15_eventsourceflex240_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s10 = irqarray15_eventsourceflex241_status;
assign irqarray15_nc_b15s11 = irqarray15_eventsourceflex241_pending;
always @(*) begin
    irqarray15_eventsourceflex241_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[1])) begin
        irqarray15_eventsourceflex241_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s20 = irqarray15_eventsourceflex242_status;
assign irqarray15_nc_b15s21 = irqarray15_eventsourceflex242_pending;
always @(*) begin
    irqarray15_eventsourceflex242_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[2])) begin
        irqarray15_eventsourceflex242_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s30 = irqarray15_eventsourceflex243_status;
assign irqarray15_nc_b15s31 = irqarray15_eventsourceflex243_pending;
always @(*) begin
    irqarray15_eventsourceflex243_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[3])) begin
        irqarray15_eventsourceflex243_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s40 = irqarray15_eventsourceflex244_status;
assign irqarray15_nc_b15s41 = irqarray15_eventsourceflex244_pending;
always @(*) begin
    irqarray15_eventsourceflex244_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[4])) begin
        irqarray15_eventsourceflex244_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s50 = irqarray15_eventsourceflex245_status;
assign irqarray15_nc_b15s51 = irqarray15_eventsourceflex245_pending;
always @(*) begin
    irqarray15_eventsourceflex245_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[5])) begin
        irqarray15_eventsourceflex245_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s60 = irqarray15_eventsourceflex246_status;
assign irqarray15_nc_b15s61 = irqarray15_eventsourceflex246_pending;
always @(*) begin
    irqarray15_eventsourceflex246_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[6])) begin
        irqarray15_eventsourceflex246_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s70 = irqarray15_eventsourceflex247_status;
assign irqarray15_nc_b15s71 = irqarray15_eventsourceflex247_pending;
always @(*) begin
    irqarray15_eventsourceflex247_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[7])) begin
        irqarray15_eventsourceflex247_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s80 = irqarray15_eventsourceflex248_status;
assign irqarray15_nc_b15s81 = irqarray15_eventsourceflex248_pending;
always @(*) begin
    irqarray15_eventsourceflex248_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[8])) begin
        irqarray15_eventsourceflex248_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s90 = irqarray15_eventsourceflex249_status;
assign irqarray15_nc_b15s91 = irqarray15_eventsourceflex249_pending;
always @(*) begin
    irqarray15_eventsourceflex249_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[9])) begin
        irqarray15_eventsourceflex249_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s100 = irqarray15_eventsourceflex250_status;
assign irqarray15_nc_b15s101 = irqarray15_eventsourceflex250_pending;
always @(*) begin
    irqarray15_eventsourceflex250_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[10])) begin
        irqarray15_eventsourceflex250_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s110 = irqarray15_eventsourceflex251_status;
assign irqarray15_nc_b15s111 = irqarray15_eventsourceflex251_pending;
always @(*) begin
    irqarray15_eventsourceflex251_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[11])) begin
        irqarray15_eventsourceflex251_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s120 = irqarray15_eventsourceflex252_status;
assign irqarray15_nc_b15s121 = irqarray15_eventsourceflex252_pending;
always @(*) begin
    irqarray15_eventsourceflex252_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[12])) begin
        irqarray15_eventsourceflex252_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s130 = irqarray15_eventsourceflex253_status;
assign irqarray15_nc_b15s131 = irqarray15_eventsourceflex253_pending;
always @(*) begin
    irqarray15_eventsourceflex253_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[13])) begin
        irqarray15_eventsourceflex253_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s140 = irqarray15_eventsourceflex254_status;
assign irqarray15_nc_b15s141 = irqarray15_eventsourceflex254_pending;
always @(*) begin
    irqarray15_eventsourceflex254_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[14])) begin
        irqarray15_eventsourceflex254_clear <= 1'd1;
    end
end
assign irqarray15_nc_b15s150 = irqarray15_eventsourceflex255_status;
assign irqarray15_nc_b15s151 = irqarray15_eventsourceflex255_pending;
always @(*) begin
    irqarray15_eventsourceflex255_clear <= 1'd0;
    if ((irqarray15_pending_re & irqarray15_pending_r[15])) begin
        irqarray15_eventsourceflex255_clear <= 1'd1;
    end
end
assign irqarray15_irq = ((((((((((((((((irqarray15_pending_status[0] & irqarray15_enable_storage[0]) | (irqarray15_pending_status[1] & irqarray15_enable_storage[1])) | (irqarray15_pending_status[2] & irqarray15_enable_storage[2])) | (irqarray15_pending_status[3] & irqarray15_enable_storage[3])) | (irqarray15_pending_status[4] & irqarray15_enable_storage[4])) | (irqarray15_pending_status[5] & irqarray15_enable_storage[5])) | (irqarray15_pending_status[6] & irqarray15_enable_storage[6])) | (irqarray15_pending_status[7] & irqarray15_enable_storage[7])) | (irqarray15_pending_status[8] & irqarray15_enable_storage[8])) | (irqarray15_pending_status[9] & irqarray15_enable_storage[9])) | (irqarray15_pending_status[10] & irqarray15_enable_storage[10])) | (irqarray15_pending_status[11] & irqarray15_enable_storage[11])) | (irqarray15_pending_status[12] & irqarray15_enable_storage[12])) | (irqarray15_pending_status[13] & irqarray15_enable_storage[13])) | (irqarray15_pending_status[14] & irqarray15_enable_storage[14])) | (irqarray15_pending_status[15] & irqarray15_enable_storage[15]));
always @(*) begin
    irqarray15_eventsourceflex240_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[0]) begin
        if (irqarray15_rising[0]) begin
            irqarray15_eventsourceflex240_trigger_filtered <= (irqarray15_interrupts[0] & (~irqarray15_eventsourceflex240_trigger_d));
        end else begin
            irqarray15_eventsourceflex240_trigger_filtered <= ((~irqarray15_interrupts[0]) & irqarray15_eventsourceflex240_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex240_trigger_filtered <= irqarray15_interrupts[0];
    end
end
assign irqarray15_eventsourceflex240_status = (irqarray15_interrupts[0] | irqarray15_trigger[0]);
always @(*) begin
    irqarray15_eventsourceflex241_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[1]) begin
        if (irqarray15_rising[1]) begin
            irqarray15_eventsourceflex241_trigger_filtered <= (irqarray15_interrupts[1] & (~irqarray15_eventsourceflex241_trigger_d));
        end else begin
            irqarray15_eventsourceflex241_trigger_filtered <= ((~irqarray15_interrupts[1]) & irqarray15_eventsourceflex241_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex241_trigger_filtered <= irqarray15_interrupts[1];
    end
end
assign irqarray15_eventsourceflex241_status = (irqarray15_interrupts[1] | irqarray15_trigger[1]);
always @(*) begin
    irqarray15_eventsourceflex242_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[2]) begin
        if (irqarray15_rising[2]) begin
            irqarray15_eventsourceflex242_trigger_filtered <= (irqarray15_interrupts[2] & (~irqarray15_eventsourceflex242_trigger_d));
        end else begin
            irqarray15_eventsourceflex242_trigger_filtered <= ((~irqarray15_interrupts[2]) & irqarray15_eventsourceflex242_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex242_trigger_filtered <= irqarray15_interrupts[2];
    end
end
assign irqarray15_eventsourceflex242_status = (irqarray15_interrupts[2] | irqarray15_trigger[2]);
always @(*) begin
    irqarray15_eventsourceflex243_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[3]) begin
        if (irqarray15_rising[3]) begin
            irqarray15_eventsourceflex243_trigger_filtered <= (irqarray15_interrupts[3] & (~irqarray15_eventsourceflex243_trigger_d));
        end else begin
            irqarray15_eventsourceflex243_trigger_filtered <= ((~irqarray15_interrupts[3]) & irqarray15_eventsourceflex243_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex243_trigger_filtered <= irqarray15_interrupts[3];
    end
end
assign irqarray15_eventsourceflex243_status = (irqarray15_interrupts[3] | irqarray15_trigger[3]);
always @(*) begin
    irqarray15_eventsourceflex244_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[4]) begin
        if (irqarray15_rising[4]) begin
            irqarray15_eventsourceflex244_trigger_filtered <= (irqarray15_interrupts[4] & (~irqarray15_eventsourceflex244_trigger_d));
        end else begin
            irqarray15_eventsourceflex244_trigger_filtered <= ((~irqarray15_interrupts[4]) & irqarray15_eventsourceflex244_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex244_trigger_filtered <= irqarray15_interrupts[4];
    end
end
assign irqarray15_eventsourceflex244_status = (irqarray15_interrupts[4] | irqarray15_trigger[4]);
always @(*) begin
    irqarray15_eventsourceflex245_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[5]) begin
        if (irqarray15_rising[5]) begin
            irqarray15_eventsourceflex245_trigger_filtered <= (irqarray15_interrupts[5] & (~irqarray15_eventsourceflex245_trigger_d));
        end else begin
            irqarray15_eventsourceflex245_trigger_filtered <= ((~irqarray15_interrupts[5]) & irqarray15_eventsourceflex245_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex245_trigger_filtered <= irqarray15_interrupts[5];
    end
end
assign irqarray15_eventsourceflex245_status = (irqarray15_interrupts[5] | irqarray15_trigger[5]);
always @(*) begin
    irqarray15_eventsourceflex246_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[6]) begin
        if (irqarray15_rising[6]) begin
            irqarray15_eventsourceflex246_trigger_filtered <= (irqarray15_interrupts[6] & (~irqarray15_eventsourceflex246_trigger_d));
        end else begin
            irqarray15_eventsourceflex246_trigger_filtered <= ((~irqarray15_interrupts[6]) & irqarray15_eventsourceflex246_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex246_trigger_filtered <= irqarray15_interrupts[6];
    end
end
assign irqarray15_eventsourceflex246_status = (irqarray15_interrupts[6] | irqarray15_trigger[6]);
always @(*) begin
    irqarray15_eventsourceflex247_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[7]) begin
        if (irqarray15_rising[7]) begin
            irqarray15_eventsourceflex247_trigger_filtered <= (irqarray15_interrupts[7] & (~irqarray15_eventsourceflex247_trigger_d));
        end else begin
            irqarray15_eventsourceflex247_trigger_filtered <= ((~irqarray15_interrupts[7]) & irqarray15_eventsourceflex247_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex247_trigger_filtered <= irqarray15_interrupts[7];
    end
end
assign irqarray15_eventsourceflex247_status = (irqarray15_interrupts[7] | irqarray15_trigger[7]);
always @(*) begin
    irqarray15_eventsourceflex248_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[8]) begin
        if (irqarray15_rising[8]) begin
            irqarray15_eventsourceflex248_trigger_filtered <= (irqarray15_interrupts[8] & (~irqarray15_eventsourceflex248_trigger_d));
        end else begin
            irqarray15_eventsourceflex248_trigger_filtered <= ((~irqarray15_interrupts[8]) & irqarray15_eventsourceflex248_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex248_trigger_filtered <= irqarray15_interrupts[8];
    end
end
assign irqarray15_eventsourceflex248_status = (irqarray15_interrupts[8] | irqarray15_trigger[8]);
always @(*) begin
    irqarray15_eventsourceflex249_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[9]) begin
        if (irqarray15_rising[9]) begin
            irqarray15_eventsourceflex249_trigger_filtered <= (irqarray15_interrupts[9] & (~irqarray15_eventsourceflex249_trigger_d));
        end else begin
            irqarray15_eventsourceflex249_trigger_filtered <= ((~irqarray15_interrupts[9]) & irqarray15_eventsourceflex249_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex249_trigger_filtered <= irqarray15_interrupts[9];
    end
end
assign irqarray15_eventsourceflex249_status = (irqarray15_interrupts[9] | irqarray15_trigger[9]);
always @(*) begin
    irqarray15_eventsourceflex250_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[10]) begin
        if (irqarray15_rising[10]) begin
            irqarray15_eventsourceflex250_trigger_filtered <= (irqarray15_interrupts[10] & (~irqarray15_eventsourceflex250_trigger_d));
        end else begin
            irqarray15_eventsourceflex250_trigger_filtered <= ((~irqarray15_interrupts[10]) & irqarray15_eventsourceflex250_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex250_trigger_filtered <= irqarray15_interrupts[10];
    end
end
assign irqarray15_eventsourceflex250_status = (irqarray15_interrupts[10] | irqarray15_trigger[10]);
always @(*) begin
    irqarray15_eventsourceflex251_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[11]) begin
        if (irqarray15_rising[11]) begin
            irqarray15_eventsourceflex251_trigger_filtered <= (irqarray15_interrupts[11] & (~irqarray15_eventsourceflex251_trigger_d));
        end else begin
            irqarray15_eventsourceflex251_trigger_filtered <= ((~irqarray15_interrupts[11]) & irqarray15_eventsourceflex251_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex251_trigger_filtered <= irqarray15_interrupts[11];
    end
end
assign irqarray15_eventsourceflex251_status = (irqarray15_interrupts[11] | irqarray15_trigger[11]);
always @(*) begin
    irqarray15_eventsourceflex252_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[12]) begin
        if (irqarray15_rising[12]) begin
            irqarray15_eventsourceflex252_trigger_filtered <= (irqarray15_interrupts[12] & (~irqarray15_eventsourceflex252_trigger_d));
        end else begin
            irqarray15_eventsourceflex252_trigger_filtered <= ((~irqarray15_interrupts[12]) & irqarray15_eventsourceflex252_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex252_trigger_filtered <= irqarray15_interrupts[12];
    end
end
assign irqarray15_eventsourceflex252_status = (irqarray15_interrupts[12] | irqarray15_trigger[12]);
always @(*) begin
    irqarray15_eventsourceflex253_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[13]) begin
        if (irqarray15_rising[13]) begin
            irqarray15_eventsourceflex253_trigger_filtered <= (irqarray15_interrupts[13] & (~irqarray15_eventsourceflex253_trigger_d));
        end else begin
            irqarray15_eventsourceflex253_trigger_filtered <= ((~irqarray15_interrupts[13]) & irqarray15_eventsourceflex253_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex253_trigger_filtered <= irqarray15_interrupts[13];
    end
end
assign irqarray15_eventsourceflex253_status = (irqarray15_interrupts[13] | irqarray15_trigger[13]);
always @(*) begin
    irqarray15_eventsourceflex254_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[14]) begin
        if (irqarray15_rising[14]) begin
            irqarray15_eventsourceflex254_trigger_filtered <= (irqarray15_interrupts[14] & (~irqarray15_eventsourceflex254_trigger_d));
        end else begin
            irqarray15_eventsourceflex254_trigger_filtered <= ((~irqarray15_interrupts[14]) & irqarray15_eventsourceflex254_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex254_trigger_filtered <= irqarray15_interrupts[14];
    end
end
assign irqarray15_eventsourceflex254_status = (irqarray15_interrupts[14] | irqarray15_trigger[14]);
always @(*) begin
    irqarray15_eventsourceflex255_trigger_filtered <= 1'd0;
    if (irqarray15_use_edge[15]) begin
        if (irqarray15_rising[15]) begin
            irqarray15_eventsourceflex255_trigger_filtered <= (irqarray15_interrupts[15] & (~irqarray15_eventsourceflex255_trigger_d));
        end else begin
            irqarray15_eventsourceflex255_trigger_filtered <= ((~irqarray15_interrupts[15]) & irqarray15_eventsourceflex255_trigger_d);
        end
    end else begin
        irqarray15_eventsourceflex255_trigger_filtered <= irqarray15_interrupts[15];
    end
end
assign irqarray15_eventsourceflex255_status = (irqarray15_interrupts[15] | irqarray15_trigger[15]);
assign irqarray16_interrupts = irq_remap16;
assign irqarray16_cam_rx_dupe0 = irqarray16_eventsourceflex256_status;
assign irqarray16_cam_rx_dupe1 = irqarray16_eventsourceflex256_pending;
always @(*) begin
    irqarray16_eventsourceflex256_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[0])) begin
        irqarray16_eventsourceflex256_clear <= 1'd1;
    end
end
assign irqarray16_i2s_rx_dupe0 = irqarray16_eventsourceflex257_status;
assign irqarray16_i2s_rx_dupe1 = irqarray16_eventsourceflex257_pending;
always @(*) begin
    irqarray16_eventsourceflex257_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[1])) begin
        irqarray16_eventsourceflex257_clear <= 1'd1;
    end
end
assign irqarray16_i2s_tx_dupe0 = irqarray16_eventsourceflex258_status;
assign irqarray16_i2s_tx_dupe1 = irqarray16_eventsourceflex258_pending;
always @(*) begin
    irqarray16_eventsourceflex258_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[2])) begin
        irqarray16_eventsourceflex258_clear <= 1'd1;
    end
end
assign irqarray16_nc_b16s30 = irqarray16_eventsourceflex259_status;
assign irqarray16_nc_b16s31 = irqarray16_eventsourceflex259_pending;
always @(*) begin
    irqarray16_eventsourceflex259_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[3])) begin
        irqarray16_eventsourceflex259_clear <= 1'd1;
    end
end
assign irqarray16_spim1_rx_dupe0 = irqarray16_eventsourceflex260_status;
assign irqarray16_spim1_rx_dupe1 = irqarray16_eventsourceflex260_pending;
always @(*) begin
    irqarray16_eventsourceflex260_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[4])) begin
        irqarray16_eventsourceflex260_clear <= 1'd1;
    end
end
assign irqarray16_spim1_tx_dupe0 = irqarray16_eventsourceflex261_status;
assign irqarray16_spim1_tx_dupe1 = irqarray16_eventsourceflex261_pending;
always @(*) begin
    irqarray16_eventsourceflex261_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[5])) begin
        irqarray16_eventsourceflex261_clear <= 1'd1;
    end
end
assign irqarray16_spim1_cmd_dupe0 = irqarray16_eventsourceflex262_status;
assign irqarray16_spim1_cmd_dupe1 = irqarray16_eventsourceflex262_pending;
always @(*) begin
    irqarray16_eventsourceflex262_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[6])) begin
        irqarray16_eventsourceflex262_clear <= 1'd1;
    end
end
assign irqarray16_spim1_eot_dupe0 = irqarray16_eventsourceflex263_status;
assign irqarray16_spim1_eot_dupe1 = irqarray16_eventsourceflex263_pending;
always @(*) begin
    irqarray16_eventsourceflex263_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[7])) begin
        irqarray16_eventsourceflex263_clear <= 1'd1;
    end
end
assign irqarray16_spim2_rx_dupe0 = irqarray16_eventsourceflex264_status;
assign irqarray16_spim2_rx_dupe1 = irqarray16_eventsourceflex264_pending;
always @(*) begin
    irqarray16_eventsourceflex264_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[8])) begin
        irqarray16_eventsourceflex264_clear <= 1'd1;
    end
end
assign irqarray16_spim2_tx_dupe0 = irqarray16_eventsourceflex265_status;
assign irqarray16_spim2_tx_dupe1 = irqarray16_eventsourceflex265_pending;
always @(*) begin
    irqarray16_eventsourceflex265_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[9])) begin
        irqarray16_eventsourceflex265_clear <= 1'd1;
    end
end
assign irqarray16_spim2_cmd_dupe0 = irqarray16_eventsourceflex266_status;
assign irqarray16_spim2_cmd_dupe1 = irqarray16_eventsourceflex266_pending;
always @(*) begin
    irqarray16_eventsourceflex266_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[10])) begin
        irqarray16_eventsourceflex266_clear <= 1'd1;
    end
end
assign irqarray16_spim2_eot_dupe0 = irqarray16_eventsourceflex267_status;
assign irqarray16_spim2_eot_dupe1 = irqarray16_eventsourceflex267_pending;
always @(*) begin
    irqarray16_eventsourceflex267_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[11])) begin
        irqarray16_eventsourceflex267_clear <= 1'd1;
    end
end
assign irqarray16_i2c0_rx_dupe0 = irqarray16_eventsourceflex268_status;
assign irqarray16_i2c0_rx_dupe1 = irqarray16_eventsourceflex268_pending;
always @(*) begin
    irqarray16_eventsourceflex268_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[12])) begin
        irqarray16_eventsourceflex268_clear <= 1'd1;
    end
end
assign irqarray16_i2c0_tx_dupe0 = irqarray16_eventsourceflex269_status;
assign irqarray16_i2c0_tx_dupe1 = irqarray16_eventsourceflex269_pending;
always @(*) begin
    irqarray16_eventsourceflex269_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[13])) begin
        irqarray16_eventsourceflex269_clear <= 1'd1;
    end
end
assign irqarray16_i2c0_cmd_dupe0 = irqarray16_eventsourceflex270_status;
assign irqarray16_i2c0_cmd_dupe1 = irqarray16_eventsourceflex270_pending;
always @(*) begin
    irqarray16_eventsourceflex270_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[14])) begin
        irqarray16_eventsourceflex270_clear <= 1'd1;
    end
end
assign irqarray16_i2c0_eot_dupe0 = irqarray16_eventsourceflex271_status;
assign irqarray16_i2c0_eot_dupe1 = irqarray16_eventsourceflex271_pending;
always @(*) begin
    irqarray16_eventsourceflex271_clear <= 1'd0;
    if ((irqarray16_pending_re & irqarray16_pending_r[15])) begin
        irqarray16_eventsourceflex271_clear <= 1'd1;
    end
end
assign irqarray16_irq = ((((((((((((((((irqarray16_pending_status[0] & irqarray16_enable_storage[0]) | (irqarray16_pending_status[1] & irqarray16_enable_storage[1])) | (irqarray16_pending_status[2] & irqarray16_enable_storage[2])) | (irqarray16_pending_status[3] & irqarray16_enable_storage[3])) | (irqarray16_pending_status[4] & irqarray16_enable_storage[4])) | (irqarray16_pending_status[5] & irqarray16_enable_storage[5])) | (irqarray16_pending_status[6] & irqarray16_enable_storage[6])) | (irqarray16_pending_status[7] & irqarray16_enable_storage[7])) | (irqarray16_pending_status[8] & irqarray16_enable_storage[8])) | (irqarray16_pending_status[9] & irqarray16_enable_storage[9])) | (irqarray16_pending_status[10] & irqarray16_enable_storage[10])) | (irqarray16_pending_status[11] & irqarray16_enable_storage[11])) | (irqarray16_pending_status[12] & irqarray16_enable_storage[12])) | (irqarray16_pending_status[13] & irqarray16_enable_storage[13])) | (irqarray16_pending_status[14] & irqarray16_enable_storage[14])) | (irqarray16_pending_status[15] & irqarray16_enable_storage[15]));
always @(*) begin
    irqarray16_eventsourceflex256_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[0]) begin
        if (irqarray16_rising[0]) begin
            irqarray16_eventsourceflex256_trigger_filtered <= (irqarray16_interrupts[0] & (~irqarray16_eventsourceflex256_trigger_d));
        end else begin
            irqarray16_eventsourceflex256_trigger_filtered <= ((~irqarray16_interrupts[0]) & irqarray16_eventsourceflex256_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex256_trigger_filtered <= irqarray16_interrupts[0];
    end
end
assign irqarray16_eventsourceflex256_status = (irqarray16_interrupts[0] | irqarray16_trigger[0]);
always @(*) begin
    irqarray16_eventsourceflex257_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[1]) begin
        if (irqarray16_rising[1]) begin
            irqarray16_eventsourceflex257_trigger_filtered <= (irqarray16_interrupts[1] & (~irqarray16_eventsourceflex257_trigger_d));
        end else begin
            irqarray16_eventsourceflex257_trigger_filtered <= ((~irqarray16_interrupts[1]) & irqarray16_eventsourceflex257_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex257_trigger_filtered <= irqarray16_interrupts[1];
    end
end
assign irqarray16_eventsourceflex257_status = (irqarray16_interrupts[1] | irqarray16_trigger[1]);
always @(*) begin
    irqarray16_eventsourceflex258_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[2]) begin
        if (irqarray16_rising[2]) begin
            irqarray16_eventsourceflex258_trigger_filtered <= (irqarray16_interrupts[2] & (~irqarray16_eventsourceflex258_trigger_d));
        end else begin
            irqarray16_eventsourceflex258_trigger_filtered <= ((~irqarray16_interrupts[2]) & irqarray16_eventsourceflex258_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex258_trigger_filtered <= irqarray16_interrupts[2];
    end
end
assign irqarray16_eventsourceflex258_status = (irqarray16_interrupts[2] | irqarray16_trigger[2]);
always @(*) begin
    irqarray16_eventsourceflex259_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[3]) begin
        if (irqarray16_rising[3]) begin
            irqarray16_eventsourceflex259_trigger_filtered <= (irqarray16_interrupts[3] & (~irqarray16_eventsourceflex259_trigger_d));
        end else begin
            irqarray16_eventsourceflex259_trigger_filtered <= ((~irqarray16_interrupts[3]) & irqarray16_eventsourceflex259_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex259_trigger_filtered <= irqarray16_interrupts[3];
    end
end
assign irqarray16_eventsourceflex259_status = (irqarray16_interrupts[3] | irqarray16_trigger[3]);
always @(*) begin
    irqarray16_eventsourceflex260_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[4]) begin
        if (irqarray16_rising[4]) begin
            irqarray16_eventsourceflex260_trigger_filtered <= (irqarray16_interrupts[4] & (~irqarray16_eventsourceflex260_trigger_d));
        end else begin
            irqarray16_eventsourceflex260_trigger_filtered <= ((~irqarray16_interrupts[4]) & irqarray16_eventsourceflex260_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex260_trigger_filtered <= irqarray16_interrupts[4];
    end
end
assign irqarray16_eventsourceflex260_status = (irqarray16_interrupts[4] | irqarray16_trigger[4]);
always @(*) begin
    irqarray16_eventsourceflex261_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[5]) begin
        if (irqarray16_rising[5]) begin
            irqarray16_eventsourceflex261_trigger_filtered <= (irqarray16_interrupts[5] & (~irqarray16_eventsourceflex261_trigger_d));
        end else begin
            irqarray16_eventsourceflex261_trigger_filtered <= ((~irqarray16_interrupts[5]) & irqarray16_eventsourceflex261_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex261_trigger_filtered <= irqarray16_interrupts[5];
    end
end
assign irqarray16_eventsourceflex261_status = (irqarray16_interrupts[5] | irqarray16_trigger[5]);
always @(*) begin
    irqarray16_eventsourceflex262_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[6]) begin
        if (irqarray16_rising[6]) begin
            irqarray16_eventsourceflex262_trigger_filtered <= (irqarray16_interrupts[6] & (~irqarray16_eventsourceflex262_trigger_d));
        end else begin
            irqarray16_eventsourceflex262_trigger_filtered <= ((~irqarray16_interrupts[6]) & irqarray16_eventsourceflex262_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex262_trigger_filtered <= irqarray16_interrupts[6];
    end
end
assign irqarray16_eventsourceflex262_status = (irqarray16_interrupts[6] | irqarray16_trigger[6]);
always @(*) begin
    irqarray16_eventsourceflex263_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[7]) begin
        if (irqarray16_rising[7]) begin
            irqarray16_eventsourceflex263_trigger_filtered <= (irqarray16_interrupts[7] & (~irqarray16_eventsourceflex263_trigger_d));
        end else begin
            irqarray16_eventsourceflex263_trigger_filtered <= ((~irqarray16_interrupts[7]) & irqarray16_eventsourceflex263_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex263_trigger_filtered <= irqarray16_interrupts[7];
    end
end
assign irqarray16_eventsourceflex263_status = (irqarray16_interrupts[7] | irqarray16_trigger[7]);
always @(*) begin
    irqarray16_eventsourceflex264_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[8]) begin
        if (irqarray16_rising[8]) begin
            irqarray16_eventsourceflex264_trigger_filtered <= (irqarray16_interrupts[8] & (~irqarray16_eventsourceflex264_trigger_d));
        end else begin
            irqarray16_eventsourceflex264_trigger_filtered <= ((~irqarray16_interrupts[8]) & irqarray16_eventsourceflex264_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex264_trigger_filtered <= irqarray16_interrupts[8];
    end
end
assign irqarray16_eventsourceflex264_status = (irqarray16_interrupts[8] | irqarray16_trigger[8]);
always @(*) begin
    irqarray16_eventsourceflex265_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[9]) begin
        if (irqarray16_rising[9]) begin
            irqarray16_eventsourceflex265_trigger_filtered <= (irqarray16_interrupts[9] & (~irqarray16_eventsourceflex265_trigger_d));
        end else begin
            irqarray16_eventsourceflex265_trigger_filtered <= ((~irqarray16_interrupts[9]) & irqarray16_eventsourceflex265_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex265_trigger_filtered <= irqarray16_interrupts[9];
    end
end
assign irqarray16_eventsourceflex265_status = (irqarray16_interrupts[9] | irqarray16_trigger[9]);
always @(*) begin
    irqarray16_eventsourceflex266_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[10]) begin
        if (irqarray16_rising[10]) begin
            irqarray16_eventsourceflex266_trigger_filtered <= (irqarray16_interrupts[10] & (~irqarray16_eventsourceflex266_trigger_d));
        end else begin
            irqarray16_eventsourceflex266_trigger_filtered <= ((~irqarray16_interrupts[10]) & irqarray16_eventsourceflex266_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex266_trigger_filtered <= irqarray16_interrupts[10];
    end
end
assign irqarray16_eventsourceflex266_status = (irqarray16_interrupts[10] | irqarray16_trigger[10]);
always @(*) begin
    irqarray16_eventsourceflex267_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[11]) begin
        if (irqarray16_rising[11]) begin
            irqarray16_eventsourceflex267_trigger_filtered <= (irqarray16_interrupts[11] & (~irqarray16_eventsourceflex267_trigger_d));
        end else begin
            irqarray16_eventsourceflex267_trigger_filtered <= ((~irqarray16_interrupts[11]) & irqarray16_eventsourceflex267_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex267_trigger_filtered <= irqarray16_interrupts[11];
    end
end
assign irqarray16_eventsourceflex267_status = (irqarray16_interrupts[11] | irqarray16_trigger[11]);
always @(*) begin
    irqarray16_eventsourceflex268_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[12]) begin
        if (irqarray16_rising[12]) begin
            irqarray16_eventsourceflex268_trigger_filtered <= (irqarray16_interrupts[12] & (~irqarray16_eventsourceflex268_trigger_d));
        end else begin
            irqarray16_eventsourceflex268_trigger_filtered <= ((~irqarray16_interrupts[12]) & irqarray16_eventsourceflex268_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex268_trigger_filtered <= irqarray16_interrupts[12];
    end
end
assign irqarray16_eventsourceflex268_status = (irqarray16_interrupts[12] | irqarray16_trigger[12]);
always @(*) begin
    irqarray16_eventsourceflex269_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[13]) begin
        if (irqarray16_rising[13]) begin
            irqarray16_eventsourceflex269_trigger_filtered <= (irqarray16_interrupts[13] & (~irqarray16_eventsourceflex269_trigger_d));
        end else begin
            irqarray16_eventsourceflex269_trigger_filtered <= ((~irqarray16_interrupts[13]) & irqarray16_eventsourceflex269_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex269_trigger_filtered <= irqarray16_interrupts[13];
    end
end
assign irqarray16_eventsourceflex269_status = (irqarray16_interrupts[13] | irqarray16_trigger[13]);
always @(*) begin
    irqarray16_eventsourceflex270_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[14]) begin
        if (irqarray16_rising[14]) begin
            irqarray16_eventsourceflex270_trigger_filtered <= (irqarray16_interrupts[14] & (~irqarray16_eventsourceflex270_trigger_d));
        end else begin
            irqarray16_eventsourceflex270_trigger_filtered <= ((~irqarray16_interrupts[14]) & irqarray16_eventsourceflex270_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex270_trigger_filtered <= irqarray16_interrupts[14];
    end
end
assign irqarray16_eventsourceflex270_status = (irqarray16_interrupts[14] | irqarray16_trigger[14]);
always @(*) begin
    irqarray16_eventsourceflex271_trigger_filtered <= 1'd0;
    if (irqarray16_use_edge[15]) begin
        if (irqarray16_rising[15]) begin
            irqarray16_eventsourceflex271_trigger_filtered <= (irqarray16_interrupts[15] & (~irqarray16_eventsourceflex271_trigger_d));
        end else begin
            irqarray16_eventsourceflex271_trigger_filtered <= ((~irqarray16_interrupts[15]) & irqarray16_eventsourceflex271_trigger_d);
        end
    end else begin
        irqarray16_eventsourceflex271_trigger_filtered <= irqarray16_interrupts[15];
    end
end
assign irqarray16_eventsourceflex271_status = (irqarray16_interrupts[15] | irqarray16_trigger[15]);
assign irqarray17_interrupts = irq_remap17;
assign irqarray17_i2c1_rx_dupe0 = irqarray17_eventsourceflex272_status;
assign irqarray17_i2c1_rx_dupe1 = irqarray17_eventsourceflex272_pending;
always @(*) begin
    irqarray17_eventsourceflex272_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[0])) begin
        irqarray17_eventsourceflex272_clear <= 1'd1;
    end
end
assign irqarray17_i2c1_tx_dupe0 = irqarray17_eventsourceflex273_status;
assign irqarray17_i2c1_tx_dupe1 = irqarray17_eventsourceflex273_pending;
always @(*) begin
    irqarray17_eventsourceflex273_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[1])) begin
        irqarray17_eventsourceflex273_clear <= 1'd1;
    end
end
assign irqarray17_i2c1_cmd_dupe0 = irqarray17_eventsourceflex274_status;
assign irqarray17_i2c1_cmd_dupe1 = irqarray17_eventsourceflex274_pending;
always @(*) begin
    irqarray17_eventsourceflex274_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[2])) begin
        irqarray17_eventsourceflex274_clear <= 1'd1;
    end
end
assign irqarray17_i2c1_eot_dupe0 = irqarray17_eventsourceflex275_status;
assign irqarray17_i2c1_eot_dupe1 = irqarray17_eventsourceflex275_pending;
always @(*) begin
    irqarray17_eventsourceflex275_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[3])) begin
        irqarray17_eventsourceflex275_clear <= 1'd1;
    end
end
assign irqarray17_pioirq0_dupe0 = irqarray17_eventsourceflex276_status;
assign irqarray17_pioirq0_dupe1 = irqarray17_eventsourceflex276_pending;
always @(*) begin
    irqarray17_eventsourceflex276_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[4])) begin
        irqarray17_eventsourceflex276_clear <= 1'd1;
    end
end
assign irqarray17_pioirq1_dupe0 = irqarray17_eventsourceflex277_status;
assign irqarray17_pioirq1_dupe1 = irqarray17_eventsourceflex277_pending;
always @(*) begin
    irqarray17_eventsourceflex277_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[5])) begin
        irqarray17_eventsourceflex277_clear <= 1'd1;
    end
end
assign irqarray17_pioirq2_dupe0 = irqarray17_eventsourceflex278_status;
assign irqarray17_pioirq2_dupe1 = irqarray17_eventsourceflex278_pending;
always @(*) begin
    irqarray17_eventsourceflex278_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[6])) begin
        irqarray17_eventsourceflex278_clear <= 1'd1;
    end
end
assign irqarray17_pioirq3_dupe0 = irqarray17_eventsourceflex279_status;
assign irqarray17_pioirq3_dupe1 = irqarray17_eventsourceflex279_pending;
always @(*) begin
    irqarray17_eventsourceflex279_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[7])) begin
        irqarray17_eventsourceflex279_clear <= 1'd1;
    end
end
assign irqarray17_qfcirq_dupe0 = irqarray17_eventsourceflex280_status;
assign irqarray17_qfcirq_dupe1 = irqarray17_eventsourceflex280_pending;
always @(*) begin
    irqarray17_eventsourceflex280_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[8])) begin
        irqarray17_eventsourceflex280_clear <= 1'd1;
    end
end
assign irqarray17_adc_rx_dupe0 = irqarray17_eventsourceflex281_status;
assign irqarray17_adc_rx_dupe1 = irqarray17_eventsourceflex281_pending;
always @(*) begin
    irqarray17_eventsourceflex281_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[9])) begin
        irqarray17_eventsourceflex281_clear <= 1'd1;
    end
end
assign irqarray17_ioxirq_dupe0 = irqarray17_eventsourceflex282_status;
assign irqarray17_ioxirq_dupe1 = irqarray17_eventsourceflex282_pending;
always @(*) begin
    irqarray17_eventsourceflex282_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[10])) begin
        irqarray17_eventsourceflex282_clear <= 1'd1;
    end
end
assign irqarray17_sddcirq_dupe0 = irqarray17_eventsourceflex283_status;
assign irqarray17_sddcirq_dupe1 = irqarray17_eventsourceflex283_pending;
always @(*) begin
    irqarray17_eventsourceflex283_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[11])) begin
        irqarray17_eventsourceflex283_clear <= 1'd1;
    end
end
assign irqarray17_nc_b17s120 = irqarray17_eventsourceflex284_status;
assign irqarray17_nc_b17s121 = irqarray17_eventsourceflex284_pending;
always @(*) begin
    irqarray17_eventsourceflex284_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[12])) begin
        irqarray17_eventsourceflex284_clear <= 1'd1;
    end
end
assign irqarray17_nc_b17s130 = irqarray17_eventsourceflex285_status;
assign irqarray17_nc_b17s131 = irqarray17_eventsourceflex285_pending;
always @(*) begin
    irqarray17_eventsourceflex285_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[13])) begin
        irqarray17_eventsourceflex285_clear <= 1'd1;
    end
end
assign irqarray17_nc_b17s140 = irqarray17_eventsourceflex286_status;
assign irqarray17_nc_b17s141 = irqarray17_eventsourceflex286_pending;
always @(*) begin
    irqarray17_eventsourceflex286_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[14])) begin
        irqarray17_eventsourceflex286_clear <= 1'd1;
    end
end
assign irqarray17_nc_b17s150 = irqarray17_eventsourceflex287_status;
assign irqarray17_nc_b17s151 = irqarray17_eventsourceflex287_pending;
always @(*) begin
    irqarray17_eventsourceflex287_clear <= 1'd0;
    if ((irqarray17_pending_re & irqarray17_pending_r[15])) begin
        irqarray17_eventsourceflex287_clear <= 1'd1;
    end
end
assign irqarray17_irq = ((((((((((((((((irqarray17_pending_status[0] & irqarray17_enable_storage[0]) | (irqarray17_pending_status[1] & irqarray17_enable_storage[1])) | (irqarray17_pending_status[2] & irqarray17_enable_storage[2])) | (irqarray17_pending_status[3] & irqarray17_enable_storage[3])) | (irqarray17_pending_status[4] & irqarray17_enable_storage[4])) | (irqarray17_pending_status[5] & irqarray17_enable_storage[5])) | (irqarray17_pending_status[6] & irqarray17_enable_storage[6])) | (irqarray17_pending_status[7] & irqarray17_enable_storage[7])) | (irqarray17_pending_status[8] & irqarray17_enable_storage[8])) | (irqarray17_pending_status[9] & irqarray17_enable_storage[9])) | (irqarray17_pending_status[10] & irqarray17_enable_storage[10])) | (irqarray17_pending_status[11] & irqarray17_enable_storage[11])) | (irqarray17_pending_status[12] & irqarray17_enable_storage[12])) | (irqarray17_pending_status[13] & irqarray17_enable_storage[13])) | (irqarray17_pending_status[14] & irqarray17_enable_storage[14])) | (irqarray17_pending_status[15] & irqarray17_enable_storage[15]));
always @(*) begin
    irqarray17_eventsourceflex272_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[0]) begin
        if (irqarray17_rising[0]) begin
            irqarray17_eventsourceflex272_trigger_filtered <= (irqarray17_interrupts[0] & (~irqarray17_eventsourceflex272_trigger_d));
        end else begin
            irqarray17_eventsourceflex272_trigger_filtered <= ((~irqarray17_interrupts[0]) & irqarray17_eventsourceflex272_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex272_trigger_filtered <= irqarray17_interrupts[0];
    end
end
assign irqarray17_eventsourceflex272_status = (irqarray17_interrupts[0] | irqarray17_trigger[0]);
always @(*) begin
    irqarray17_eventsourceflex273_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[1]) begin
        if (irqarray17_rising[1]) begin
            irqarray17_eventsourceflex273_trigger_filtered <= (irqarray17_interrupts[1] & (~irqarray17_eventsourceflex273_trigger_d));
        end else begin
            irqarray17_eventsourceflex273_trigger_filtered <= ((~irqarray17_interrupts[1]) & irqarray17_eventsourceflex273_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex273_trigger_filtered <= irqarray17_interrupts[1];
    end
end
assign irqarray17_eventsourceflex273_status = (irqarray17_interrupts[1] | irqarray17_trigger[1]);
always @(*) begin
    irqarray17_eventsourceflex274_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[2]) begin
        if (irqarray17_rising[2]) begin
            irqarray17_eventsourceflex274_trigger_filtered <= (irqarray17_interrupts[2] & (~irqarray17_eventsourceflex274_trigger_d));
        end else begin
            irqarray17_eventsourceflex274_trigger_filtered <= ((~irqarray17_interrupts[2]) & irqarray17_eventsourceflex274_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex274_trigger_filtered <= irqarray17_interrupts[2];
    end
end
assign irqarray17_eventsourceflex274_status = (irqarray17_interrupts[2] | irqarray17_trigger[2]);
always @(*) begin
    irqarray17_eventsourceflex275_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[3]) begin
        if (irqarray17_rising[3]) begin
            irqarray17_eventsourceflex275_trigger_filtered <= (irqarray17_interrupts[3] & (~irqarray17_eventsourceflex275_trigger_d));
        end else begin
            irqarray17_eventsourceflex275_trigger_filtered <= ((~irqarray17_interrupts[3]) & irqarray17_eventsourceflex275_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex275_trigger_filtered <= irqarray17_interrupts[3];
    end
end
assign irqarray17_eventsourceflex275_status = (irqarray17_interrupts[3] | irqarray17_trigger[3]);
always @(*) begin
    irqarray17_eventsourceflex276_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[4]) begin
        if (irqarray17_rising[4]) begin
            irqarray17_eventsourceflex276_trigger_filtered <= (irqarray17_interrupts[4] & (~irqarray17_eventsourceflex276_trigger_d));
        end else begin
            irqarray17_eventsourceflex276_trigger_filtered <= ((~irqarray17_interrupts[4]) & irqarray17_eventsourceflex276_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex276_trigger_filtered <= irqarray17_interrupts[4];
    end
end
assign irqarray17_eventsourceflex276_status = (irqarray17_interrupts[4] | irqarray17_trigger[4]);
always @(*) begin
    irqarray17_eventsourceflex277_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[5]) begin
        if (irqarray17_rising[5]) begin
            irqarray17_eventsourceflex277_trigger_filtered <= (irqarray17_interrupts[5] & (~irqarray17_eventsourceflex277_trigger_d));
        end else begin
            irqarray17_eventsourceflex277_trigger_filtered <= ((~irqarray17_interrupts[5]) & irqarray17_eventsourceflex277_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex277_trigger_filtered <= irqarray17_interrupts[5];
    end
end
assign irqarray17_eventsourceflex277_status = (irqarray17_interrupts[5] | irqarray17_trigger[5]);
always @(*) begin
    irqarray17_eventsourceflex278_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[6]) begin
        if (irqarray17_rising[6]) begin
            irqarray17_eventsourceflex278_trigger_filtered <= (irqarray17_interrupts[6] & (~irqarray17_eventsourceflex278_trigger_d));
        end else begin
            irqarray17_eventsourceflex278_trigger_filtered <= ((~irqarray17_interrupts[6]) & irqarray17_eventsourceflex278_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex278_trigger_filtered <= irqarray17_interrupts[6];
    end
end
assign irqarray17_eventsourceflex278_status = (irqarray17_interrupts[6] | irqarray17_trigger[6]);
always @(*) begin
    irqarray17_eventsourceflex279_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[7]) begin
        if (irqarray17_rising[7]) begin
            irqarray17_eventsourceflex279_trigger_filtered <= (irqarray17_interrupts[7] & (~irqarray17_eventsourceflex279_trigger_d));
        end else begin
            irqarray17_eventsourceflex279_trigger_filtered <= ((~irqarray17_interrupts[7]) & irqarray17_eventsourceflex279_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex279_trigger_filtered <= irqarray17_interrupts[7];
    end
end
assign irqarray17_eventsourceflex279_status = (irqarray17_interrupts[7] | irqarray17_trigger[7]);
always @(*) begin
    irqarray17_eventsourceflex280_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[8]) begin
        if (irqarray17_rising[8]) begin
            irqarray17_eventsourceflex280_trigger_filtered <= (irqarray17_interrupts[8] & (~irqarray17_eventsourceflex280_trigger_d));
        end else begin
            irqarray17_eventsourceflex280_trigger_filtered <= ((~irqarray17_interrupts[8]) & irqarray17_eventsourceflex280_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex280_trigger_filtered <= irqarray17_interrupts[8];
    end
end
assign irqarray17_eventsourceflex280_status = (irqarray17_interrupts[8] | irqarray17_trigger[8]);
always @(*) begin
    irqarray17_eventsourceflex281_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[9]) begin
        if (irqarray17_rising[9]) begin
            irqarray17_eventsourceflex281_trigger_filtered <= (irqarray17_interrupts[9] & (~irqarray17_eventsourceflex281_trigger_d));
        end else begin
            irqarray17_eventsourceflex281_trigger_filtered <= ((~irqarray17_interrupts[9]) & irqarray17_eventsourceflex281_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex281_trigger_filtered <= irqarray17_interrupts[9];
    end
end
assign irqarray17_eventsourceflex281_status = (irqarray17_interrupts[9] | irqarray17_trigger[9]);
always @(*) begin
    irqarray17_eventsourceflex282_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[10]) begin
        if (irqarray17_rising[10]) begin
            irqarray17_eventsourceflex282_trigger_filtered <= (irqarray17_interrupts[10] & (~irqarray17_eventsourceflex282_trigger_d));
        end else begin
            irqarray17_eventsourceflex282_trigger_filtered <= ((~irqarray17_interrupts[10]) & irqarray17_eventsourceflex282_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex282_trigger_filtered <= irqarray17_interrupts[10];
    end
end
assign irqarray17_eventsourceflex282_status = (irqarray17_interrupts[10] | irqarray17_trigger[10]);
always @(*) begin
    irqarray17_eventsourceflex283_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[11]) begin
        if (irqarray17_rising[11]) begin
            irqarray17_eventsourceflex283_trigger_filtered <= (irqarray17_interrupts[11] & (~irqarray17_eventsourceflex283_trigger_d));
        end else begin
            irqarray17_eventsourceflex283_trigger_filtered <= ((~irqarray17_interrupts[11]) & irqarray17_eventsourceflex283_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex283_trigger_filtered <= irqarray17_interrupts[11];
    end
end
assign irqarray17_eventsourceflex283_status = (irqarray17_interrupts[11] | irqarray17_trigger[11]);
always @(*) begin
    irqarray17_eventsourceflex284_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[12]) begin
        if (irqarray17_rising[12]) begin
            irqarray17_eventsourceflex284_trigger_filtered <= (irqarray17_interrupts[12] & (~irqarray17_eventsourceflex284_trigger_d));
        end else begin
            irqarray17_eventsourceflex284_trigger_filtered <= ((~irqarray17_interrupts[12]) & irqarray17_eventsourceflex284_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex284_trigger_filtered <= irqarray17_interrupts[12];
    end
end
assign irqarray17_eventsourceflex284_status = (irqarray17_interrupts[12] | irqarray17_trigger[12]);
always @(*) begin
    irqarray17_eventsourceflex285_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[13]) begin
        if (irqarray17_rising[13]) begin
            irqarray17_eventsourceflex285_trigger_filtered <= (irqarray17_interrupts[13] & (~irqarray17_eventsourceflex285_trigger_d));
        end else begin
            irqarray17_eventsourceflex285_trigger_filtered <= ((~irqarray17_interrupts[13]) & irqarray17_eventsourceflex285_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex285_trigger_filtered <= irqarray17_interrupts[13];
    end
end
assign irqarray17_eventsourceflex285_status = (irqarray17_interrupts[13] | irqarray17_trigger[13]);
always @(*) begin
    irqarray17_eventsourceflex286_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[14]) begin
        if (irqarray17_rising[14]) begin
            irqarray17_eventsourceflex286_trigger_filtered <= (irqarray17_interrupts[14] & (~irqarray17_eventsourceflex286_trigger_d));
        end else begin
            irqarray17_eventsourceflex286_trigger_filtered <= ((~irqarray17_interrupts[14]) & irqarray17_eventsourceflex286_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex286_trigger_filtered <= irqarray17_interrupts[14];
    end
end
assign irqarray17_eventsourceflex286_status = (irqarray17_interrupts[14] | irqarray17_trigger[14]);
always @(*) begin
    irqarray17_eventsourceflex287_trigger_filtered <= 1'd0;
    if (irqarray17_use_edge[15]) begin
        if (irqarray17_rising[15]) begin
            irqarray17_eventsourceflex287_trigger_filtered <= (irqarray17_interrupts[15] & (~irqarray17_eventsourceflex287_trigger_d));
        end else begin
            irqarray17_eventsourceflex287_trigger_filtered <= ((~irqarray17_interrupts[15]) & irqarray17_eventsourceflex287_trigger_d);
        end
    end else begin
        irqarray17_eventsourceflex287_trigger_filtered <= irqarray17_interrupts[15];
    end
end
assign irqarray17_eventsourceflex287_status = (irqarray17_interrupts[15] | irqarray17_trigger[15]);
assign irqarray18_interrupts = irq_remap18;
assign irqarray18_pioirq0_dupe0 = irqarray18_eventsourceflex288_status;
assign irqarray18_pioirq0_dupe1 = irqarray18_eventsourceflex288_pending;
always @(*) begin
    irqarray18_eventsourceflex288_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[0])) begin
        irqarray18_eventsourceflex288_clear <= 1'd1;
    end
end
assign irqarray18_pioirq1_dupe0 = irqarray18_eventsourceflex289_status;
assign irqarray18_pioirq1_dupe1 = irqarray18_eventsourceflex289_pending;
always @(*) begin
    irqarray18_eventsourceflex289_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[1])) begin
        irqarray18_eventsourceflex289_clear <= 1'd1;
    end
end
assign irqarray18_pioirq2_dupe0 = irqarray18_eventsourceflex290_status;
assign irqarray18_pioirq2_dupe1 = irqarray18_eventsourceflex290_pending;
always @(*) begin
    irqarray18_eventsourceflex290_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[2])) begin
        irqarray18_eventsourceflex290_clear <= 1'd1;
    end
end
assign irqarray18_pioirq3_dupe0 = irqarray18_eventsourceflex291_status;
assign irqarray18_pioirq3_dupe1 = irqarray18_eventsourceflex291_pending;
always @(*) begin
    irqarray18_eventsourceflex291_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[3])) begin
        irqarray18_eventsourceflex291_clear <= 1'd1;
    end
end
assign irqarray18_i2c2_rx_dupe0 = irqarray18_eventsourceflex292_status;
assign irqarray18_i2c2_rx_dupe1 = irqarray18_eventsourceflex292_pending;
always @(*) begin
    irqarray18_eventsourceflex292_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[4])) begin
        irqarray18_eventsourceflex292_clear <= 1'd1;
    end
end
assign irqarray18_i2c2_tx_dupe0 = irqarray18_eventsourceflex293_status;
assign irqarray18_i2c2_tx_dupe1 = irqarray18_eventsourceflex293_pending;
always @(*) begin
    irqarray18_eventsourceflex293_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[5])) begin
        irqarray18_eventsourceflex293_clear <= 1'd1;
    end
end
assign irqarray18_i2c2_cmd_dupe0 = irqarray18_eventsourceflex294_status;
assign irqarray18_i2c2_cmd_dupe1 = irqarray18_eventsourceflex294_pending;
always @(*) begin
    irqarray18_eventsourceflex294_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[6])) begin
        irqarray18_eventsourceflex294_clear <= 1'd1;
    end
end
assign irqarray18_i2c2_eot_dupe0 = irqarray18_eventsourceflex295_status;
assign irqarray18_i2c2_eot_dupe1 = irqarray18_eventsourceflex295_pending;
always @(*) begin
    irqarray18_eventsourceflex295_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[7])) begin
        irqarray18_eventsourceflex295_clear <= 1'd1;
    end
end
assign irqarray18_i2c0_nack_dupe0 = irqarray18_eventsourceflex296_status;
assign irqarray18_i2c0_nack_dupe1 = irqarray18_eventsourceflex296_pending;
always @(*) begin
    irqarray18_eventsourceflex296_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[8])) begin
        irqarray18_eventsourceflex296_clear <= 1'd1;
    end
end
assign irqarray18_i2c1_nack_dupe0 = irqarray18_eventsourceflex297_status;
assign irqarray18_i2c1_nack_dupe1 = irqarray18_eventsourceflex297_pending;
always @(*) begin
    irqarray18_eventsourceflex297_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[9])) begin
        irqarray18_eventsourceflex297_clear <= 1'd1;
    end
end
assign irqarray18_i2c2_nack_dupe0 = irqarray18_eventsourceflex298_status;
assign irqarray18_i2c2_nack_dupe1 = irqarray18_eventsourceflex298_pending;
always @(*) begin
    irqarray18_eventsourceflex298_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[10])) begin
        irqarray18_eventsourceflex298_clear <= 1'd1;
    end
end
assign irqarray18_i2c0_err_dupe0 = irqarray18_eventsourceflex299_status;
assign irqarray18_i2c0_err_dupe1 = irqarray18_eventsourceflex299_pending;
always @(*) begin
    irqarray18_eventsourceflex299_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[11])) begin
        irqarray18_eventsourceflex299_clear <= 1'd1;
    end
end
assign irqarray18_i2c1_err_dupe0 = irqarray18_eventsourceflex300_status;
assign irqarray18_i2c1_err_dupe1 = irqarray18_eventsourceflex300_pending;
always @(*) begin
    irqarray18_eventsourceflex300_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[12])) begin
        irqarray18_eventsourceflex300_clear <= 1'd1;
    end
end
assign irqarray18_i2c2_err_dupe0 = irqarray18_eventsourceflex301_status;
assign irqarray18_i2c2_err_dupe1 = irqarray18_eventsourceflex301_pending;
always @(*) begin
    irqarray18_eventsourceflex301_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[13])) begin
        irqarray18_eventsourceflex301_clear <= 1'd1;
    end
end
assign irqarray18_ioxirq_dupe0 = irqarray18_eventsourceflex302_status;
assign irqarray18_ioxirq_dupe1 = irqarray18_eventsourceflex302_pending;
always @(*) begin
    irqarray18_eventsourceflex302_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[14])) begin
        irqarray18_eventsourceflex302_clear <= 1'd1;
    end
end
assign irqarray18_cam_rx_dupe0 = irqarray18_eventsourceflex303_status;
assign irqarray18_cam_rx_dupe1 = irqarray18_eventsourceflex303_pending;
always @(*) begin
    irqarray18_eventsourceflex303_clear <= 1'd0;
    if ((irqarray18_pending_re & irqarray18_pending_r[15])) begin
        irqarray18_eventsourceflex303_clear <= 1'd1;
    end
end
assign irqarray18_irq = ((((((((((((((((irqarray18_pending_status[0] & irqarray18_enable_storage[0]) | (irqarray18_pending_status[1] & irqarray18_enable_storage[1])) | (irqarray18_pending_status[2] & irqarray18_enable_storage[2])) | (irqarray18_pending_status[3] & irqarray18_enable_storage[3])) | (irqarray18_pending_status[4] & irqarray18_enable_storage[4])) | (irqarray18_pending_status[5] & irqarray18_enable_storage[5])) | (irqarray18_pending_status[6] & irqarray18_enable_storage[6])) | (irqarray18_pending_status[7] & irqarray18_enable_storage[7])) | (irqarray18_pending_status[8] & irqarray18_enable_storage[8])) | (irqarray18_pending_status[9] & irqarray18_enable_storage[9])) | (irqarray18_pending_status[10] & irqarray18_enable_storage[10])) | (irqarray18_pending_status[11] & irqarray18_enable_storage[11])) | (irqarray18_pending_status[12] & irqarray18_enable_storage[12])) | (irqarray18_pending_status[13] & irqarray18_enable_storage[13])) | (irqarray18_pending_status[14] & irqarray18_enable_storage[14])) | (irqarray18_pending_status[15] & irqarray18_enable_storage[15]));
always @(*) begin
    irqarray18_eventsourceflex288_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[0]) begin
        if (irqarray18_rising[0]) begin
            irqarray18_eventsourceflex288_trigger_filtered <= (irqarray18_interrupts[0] & (~irqarray18_eventsourceflex288_trigger_d));
        end else begin
            irqarray18_eventsourceflex288_trigger_filtered <= ((~irqarray18_interrupts[0]) & irqarray18_eventsourceflex288_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex288_trigger_filtered <= irqarray18_interrupts[0];
    end
end
assign irqarray18_eventsourceflex288_status = (irqarray18_interrupts[0] | irqarray18_trigger[0]);
always @(*) begin
    irqarray18_eventsourceflex289_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[1]) begin
        if (irqarray18_rising[1]) begin
            irqarray18_eventsourceflex289_trigger_filtered <= (irqarray18_interrupts[1] & (~irqarray18_eventsourceflex289_trigger_d));
        end else begin
            irqarray18_eventsourceflex289_trigger_filtered <= ((~irqarray18_interrupts[1]) & irqarray18_eventsourceflex289_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex289_trigger_filtered <= irqarray18_interrupts[1];
    end
end
assign irqarray18_eventsourceflex289_status = (irqarray18_interrupts[1] | irqarray18_trigger[1]);
always @(*) begin
    irqarray18_eventsourceflex290_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[2]) begin
        if (irqarray18_rising[2]) begin
            irqarray18_eventsourceflex290_trigger_filtered <= (irqarray18_interrupts[2] & (~irqarray18_eventsourceflex290_trigger_d));
        end else begin
            irqarray18_eventsourceflex290_trigger_filtered <= ((~irqarray18_interrupts[2]) & irqarray18_eventsourceflex290_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex290_trigger_filtered <= irqarray18_interrupts[2];
    end
end
assign irqarray18_eventsourceflex290_status = (irqarray18_interrupts[2] | irqarray18_trigger[2]);
always @(*) begin
    irqarray18_eventsourceflex291_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[3]) begin
        if (irqarray18_rising[3]) begin
            irqarray18_eventsourceflex291_trigger_filtered <= (irqarray18_interrupts[3] & (~irqarray18_eventsourceflex291_trigger_d));
        end else begin
            irqarray18_eventsourceflex291_trigger_filtered <= ((~irqarray18_interrupts[3]) & irqarray18_eventsourceflex291_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex291_trigger_filtered <= irqarray18_interrupts[3];
    end
end
assign irqarray18_eventsourceflex291_status = (irqarray18_interrupts[3] | irqarray18_trigger[3]);
always @(*) begin
    irqarray18_eventsourceflex292_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[4]) begin
        if (irqarray18_rising[4]) begin
            irqarray18_eventsourceflex292_trigger_filtered <= (irqarray18_interrupts[4] & (~irqarray18_eventsourceflex292_trigger_d));
        end else begin
            irqarray18_eventsourceflex292_trigger_filtered <= ((~irqarray18_interrupts[4]) & irqarray18_eventsourceflex292_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex292_trigger_filtered <= irqarray18_interrupts[4];
    end
end
assign irqarray18_eventsourceflex292_status = (irqarray18_interrupts[4] | irqarray18_trigger[4]);
always @(*) begin
    irqarray18_eventsourceflex293_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[5]) begin
        if (irqarray18_rising[5]) begin
            irqarray18_eventsourceflex293_trigger_filtered <= (irqarray18_interrupts[5] & (~irqarray18_eventsourceflex293_trigger_d));
        end else begin
            irqarray18_eventsourceflex293_trigger_filtered <= ((~irqarray18_interrupts[5]) & irqarray18_eventsourceflex293_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex293_trigger_filtered <= irqarray18_interrupts[5];
    end
end
assign irqarray18_eventsourceflex293_status = (irqarray18_interrupts[5] | irqarray18_trigger[5]);
always @(*) begin
    irqarray18_eventsourceflex294_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[6]) begin
        if (irqarray18_rising[6]) begin
            irqarray18_eventsourceflex294_trigger_filtered <= (irqarray18_interrupts[6] & (~irqarray18_eventsourceflex294_trigger_d));
        end else begin
            irqarray18_eventsourceflex294_trigger_filtered <= ((~irqarray18_interrupts[6]) & irqarray18_eventsourceflex294_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex294_trigger_filtered <= irqarray18_interrupts[6];
    end
end
assign irqarray18_eventsourceflex294_status = (irqarray18_interrupts[6] | irqarray18_trigger[6]);
always @(*) begin
    irqarray18_eventsourceflex295_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[7]) begin
        if (irqarray18_rising[7]) begin
            irqarray18_eventsourceflex295_trigger_filtered <= (irqarray18_interrupts[7] & (~irqarray18_eventsourceflex295_trigger_d));
        end else begin
            irqarray18_eventsourceflex295_trigger_filtered <= ((~irqarray18_interrupts[7]) & irqarray18_eventsourceflex295_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex295_trigger_filtered <= irqarray18_interrupts[7];
    end
end
assign irqarray18_eventsourceflex295_status = (irqarray18_interrupts[7] | irqarray18_trigger[7]);
always @(*) begin
    irqarray18_eventsourceflex296_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[8]) begin
        if (irqarray18_rising[8]) begin
            irqarray18_eventsourceflex296_trigger_filtered <= (irqarray18_interrupts[8] & (~irqarray18_eventsourceflex296_trigger_d));
        end else begin
            irqarray18_eventsourceflex296_trigger_filtered <= ((~irqarray18_interrupts[8]) & irqarray18_eventsourceflex296_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex296_trigger_filtered <= irqarray18_interrupts[8];
    end
end
assign irqarray18_eventsourceflex296_status = (irqarray18_interrupts[8] | irqarray18_trigger[8]);
always @(*) begin
    irqarray18_eventsourceflex297_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[9]) begin
        if (irqarray18_rising[9]) begin
            irqarray18_eventsourceflex297_trigger_filtered <= (irqarray18_interrupts[9] & (~irqarray18_eventsourceflex297_trigger_d));
        end else begin
            irqarray18_eventsourceflex297_trigger_filtered <= ((~irqarray18_interrupts[9]) & irqarray18_eventsourceflex297_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex297_trigger_filtered <= irqarray18_interrupts[9];
    end
end
assign irqarray18_eventsourceflex297_status = (irqarray18_interrupts[9] | irqarray18_trigger[9]);
always @(*) begin
    irqarray18_eventsourceflex298_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[10]) begin
        if (irqarray18_rising[10]) begin
            irqarray18_eventsourceflex298_trigger_filtered <= (irqarray18_interrupts[10] & (~irqarray18_eventsourceflex298_trigger_d));
        end else begin
            irqarray18_eventsourceflex298_trigger_filtered <= ((~irqarray18_interrupts[10]) & irqarray18_eventsourceflex298_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex298_trigger_filtered <= irqarray18_interrupts[10];
    end
end
assign irqarray18_eventsourceflex298_status = (irqarray18_interrupts[10] | irqarray18_trigger[10]);
always @(*) begin
    irqarray18_eventsourceflex299_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[11]) begin
        if (irqarray18_rising[11]) begin
            irqarray18_eventsourceflex299_trigger_filtered <= (irqarray18_interrupts[11] & (~irqarray18_eventsourceflex299_trigger_d));
        end else begin
            irqarray18_eventsourceflex299_trigger_filtered <= ((~irqarray18_interrupts[11]) & irqarray18_eventsourceflex299_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex299_trigger_filtered <= irqarray18_interrupts[11];
    end
end
assign irqarray18_eventsourceflex299_status = (irqarray18_interrupts[11] | irqarray18_trigger[11]);
always @(*) begin
    irqarray18_eventsourceflex300_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[12]) begin
        if (irqarray18_rising[12]) begin
            irqarray18_eventsourceflex300_trigger_filtered <= (irqarray18_interrupts[12] & (~irqarray18_eventsourceflex300_trigger_d));
        end else begin
            irqarray18_eventsourceflex300_trigger_filtered <= ((~irqarray18_interrupts[12]) & irqarray18_eventsourceflex300_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex300_trigger_filtered <= irqarray18_interrupts[12];
    end
end
assign irqarray18_eventsourceflex300_status = (irqarray18_interrupts[12] | irqarray18_trigger[12]);
always @(*) begin
    irqarray18_eventsourceflex301_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[13]) begin
        if (irqarray18_rising[13]) begin
            irqarray18_eventsourceflex301_trigger_filtered <= (irqarray18_interrupts[13] & (~irqarray18_eventsourceflex301_trigger_d));
        end else begin
            irqarray18_eventsourceflex301_trigger_filtered <= ((~irqarray18_interrupts[13]) & irqarray18_eventsourceflex301_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex301_trigger_filtered <= irqarray18_interrupts[13];
    end
end
assign irqarray18_eventsourceflex301_status = (irqarray18_interrupts[13] | irqarray18_trigger[13]);
always @(*) begin
    irqarray18_eventsourceflex302_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[14]) begin
        if (irqarray18_rising[14]) begin
            irqarray18_eventsourceflex302_trigger_filtered <= (irqarray18_interrupts[14] & (~irqarray18_eventsourceflex302_trigger_d));
        end else begin
            irqarray18_eventsourceflex302_trigger_filtered <= ((~irqarray18_interrupts[14]) & irqarray18_eventsourceflex302_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex302_trigger_filtered <= irqarray18_interrupts[14];
    end
end
assign irqarray18_eventsourceflex302_status = (irqarray18_interrupts[14] | irqarray18_trigger[14]);
always @(*) begin
    irqarray18_eventsourceflex303_trigger_filtered <= 1'd0;
    if (irqarray18_use_edge[15]) begin
        if (irqarray18_rising[15]) begin
            irqarray18_eventsourceflex303_trigger_filtered <= (irqarray18_interrupts[15] & (~irqarray18_eventsourceflex303_trigger_d));
        end else begin
            irqarray18_eventsourceflex303_trigger_filtered <= ((~irqarray18_interrupts[15]) & irqarray18_eventsourceflex303_trigger_d);
        end
    end else begin
        irqarray18_eventsourceflex303_trigger_filtered <= irqarray18_interrupts[15];
    end
end
assign irqarray18_eventsourceflex303_status = (irqarray18_interrupts[15] | irqarray18_trigger[15]);
assign irqarray19_interrupts = irq_remap19;
assign irqarray19_mbox_irq_available_dupe0 = irqarray19_eventsourceflex304_status;
assign irqarray19_mbox_irq_available_dupe1 = irqarray19_eventsourceflex304_pending;
always @(*) begin
    irqarray19_eventsourceflex304_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[0])) begin
        irqarray19_eventsourceflex304_clear <= 1'd1;
    end
end
assign irqarray19_mbox_irq_abort_init_dupe0 = irqarray19_eventsourceflex305_status;
assign irqarray19_mbox_irq_abort_init_dupe1 = irqarray19_eventsourceflex305_pending;
always @(*) begin
    irqarray19_eventsourceflex305_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[1])) begin
        irqarray19_eventsourceflex305_clear <= 1'd1;
    end
end
assign irqarray19_mbox_irq_done_dupe0 = irqarray19_eventsourceflex306_status;
assign irqarray19_mbox_irq_done_dupe1 = irqarray19_eventsourceflex306_pending;
always @(*) begin
    irqarray19_eventsourceflex306_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[2])) begin
        irqarray19_eventsourceflex306_clear <= 1'd1;
    end
end
assign irqarray19_mbox_irq_error_dupe0 = irqarray19_eventsourceflex307_status;
assign irqarray19_mbox_irq_error_dupe1 = irqarray19_eventsourceflex307_pending;
always @(*) begin
    irqarray19_eventsourceflex307_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[3])) begin
        irqarray19_eventsourceflex307_clear <= 1'd1;
    end
end
assign irqarray19_pioirq0_dupe0 = irqarray19_eventsourceflex308_status;
assign irqarray19_pioirq0_dupe1 = irqarray19_eventsourceflex308_pending;
always @(*) begin
    irqarray19_eventsourceflex308_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[4])) begin
        irqarray19_eventsourceflex308_clear <= 1'd1;
    end
end
assign irqarray19_pioirq1_dupe0 = irqarray19_eventsourceflex309_status;
assign irqarray19_pioirq1_dupe1 = irqarray19_eventsourceflex309_pending;
always @(*) begin
    irqarray19_eventsourceflex309_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[5])) begin
        irqarray19_eventsourceflex309_clear <= 1'd1;
    end
end
assign irqarray19_pioirq2_dupe0 = irqarray19_eventsourceflex310_status;
assign irqarray19_pioirq2_dupe1 = irqarray19_eventsourceflex310_pending;
always @(*) begin
    irqarray19_eventsourceflex310_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[6])) begin
        irqarray19_eventsourceflex310_clear <= 1'd1;
    end
end
assign irqarray19_pioirq3_dupe0 = irqarray19_eventsourceflex311_status;
assign irqarray19_pioirq3_dupe1 = irqarray19_eventsourceflex311_pending;
always @(*) begin
    irqarray19_eventsourceflex311_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[7])) begin
        irqarray19_eventsourceflex311_clear <= 1'd1;
    end
end
assign irqarray19_sdio_rx_dupe0 = irqarray19_eventsourceflex312_status;
assign irqarray19_sdio_rx_dupe1 = irqarray19_eventsourceflex312_pending;
always @(*) begin
    irqarray19_eventsourceflex312_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[8])) begin
        irqarray19_eventsourceflex312_clear <= 1'd1;
    end
end
assign irqarray19_sdio_tx_dupe0 = irqarray19_eventsourceflex313_status;
assign irqarray19_sdio_tx_dupe1 = irqarray19_eventsourceflex313_pending;
always @(*) begin
    irqarray19_eventsourceflex313_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[9])) begin
        irqarray19_eventsourceflex313_clear <= 1'd1;
    end
end
assign irqarray19_sdio_eot_dupe0 = irqarray19_eventsourceflex314_status;
assign irqarray19_sdio_eot_dupe1 = irqarray19_eventsourceflex314_pending;
always @(*) begin
    irqarray19_eventsourceflex314_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[10])) begin
        irqarray19_eventsourceflex314_clear <= 1'd1;
    end
end
assign irqarray19_sdio_err_dupe0 = irqarray19_eventsourceflex315_status;
assign irqarray19_sdio_err_dupe1 = irqarray19_eventsourceflex315_pending;
always @(*) begin
    irqarray19_eventsourceflex315_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[11])) begin
        irqarray19_eventsourceflex315_clear <= 1'd1;
    end
end
assign irqarray19_nc_b19s120 = irqarray19_eventsourceflex316_status;
assign irqarray19_nc_b19s121 = irqarray19_eventsourceflex316_pending;
always @(*) begin
    irqarray19_eventsourceflex316_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[12])) begin
        irqarray19_eventsourceflex316_clear <= 1'd1;
    end
end
assign irqarray19_nc_b19s130 = irqarray19_eventsourceflex317_status;
assign irqarray19_nc_b19s131 = irqarray19_eventsourceflex317_pending;
always @(*) begin
    irqarray19_eventsourceflex317_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[13])) begin
        irqarray19_eventsourceflex317_clear <= 1'd1;
    end
end
assign irqarray19_nc_b19s140 = irqarray19_eventsourceflex318_status;
assign irqarray19_nc_b19s141 = irqarray19_eventsourceflex318_pending;
always @(*) begin
    irqarray19_eventsourceflex318_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[14])) begin
        irqarray19_eventsourceflex318_clear <= 1'd1;
    end
end
assign irqarray19_nc_b19s150 = irqarray19_eventsourceflex319_status;
assign irqarray19_nc_b19s151 = irqarray19_eventsourceflex319_pending;
always @(*) begin
    irqarray19_eventsourceflex319_clear <= 1'd0;
    if ((irqarray19_pending_re & irqarray19_pending_r[15])) begin
        irqarray19_eventsourceflex319_clear <= 1'd1;
    end
end
assign irqarray19_irq = ((((((((((((((((irqarray19_pending_status[0] & irqarray19_enable_storage[0]) | (irqarray19_pending_status[1] & irqarray19_enable_storage[1])) | (irqarray19_pending_status[2] & irqarray19_enable_storage[2])) | (irqarray19_pending_status[3] & irqarray19_enable_storage[3])) | (irqarray19_pending_status[4] & irqarray19_enable_storage[4])) | (irqarray19_pending_status[5] & irqarray19_enable_storage[5])) | (irqarray19_pending_status[6] & irqarray19_enable_storage[6])) | (irqarray19_pending_status[7] & irqarray19_enable_storage[7])) | (irqarray19_pending_status[8] & irqarray19_enable_storage[8])) | (irqarray19_pending_status[9] & irqarray19_enable_storage[9])) | (irqarray19_pending_status[10] & irqarray19_enable_storage[10])) | (irqarray19_pending_status[11] & irqarray19_enable_storage[11])) | (irqarray19_pending_status[12] & irqarray19_enable_storage[12])) | (irqarray19_pending_status[13] & irqarray19_enable_storage[13])) | (irqarray19_pending_status[14] & irqarray19_enable_storage[14])) | (irqarray19_pending_status[15] & irqarray19_enable_storage[15]));
always @(*) begin
    irqarray19_eventsourceflex304_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[0]) begin
        if (irqarray19_rising[0]) begin
            irqarray19_eventsourceflex304_trigger_filtered <= (irqarray19_interrupts[0] & (~irqarray19_eventsourceflex304_trigger_d));
        end else begin
            irqarray19_eventsourceflex304_trigger_filtered <= ((~irqarray19_interrupts[0]) & irqarray19_eventsourceflex304_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex304_trigger_filtered <= irqarray19_interrupts[0];
    end
end
assign irqarray19_eventsourceflex304_status = (irqarray19_interrupts[0] | irqarray19_trigger[0]);
always @(*) begin
    irqarray19_eventsourceflex305_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[1]) begin
        if (irqarray19_rising[1]) begin
            irqarray19_eventsourceflex305_trigger_filtered <= (irqarray19_interrupts[1] & (~irqarray19_eventsourceflex305_trigger_d));
        end else begin
            irqarray19_eventsourceflex305_trigger_filtered <= ((~irqarray19_interrupts[1]) & irqarray19_eventsourceflex305_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex305_trigger_filtered <= irqarray19_interrupts[1];
    end
end
assign irqarray19_eventsourceflex305_status = (irqarray19_interrupts[1] | irqarray19_trigger[1]);
always @(*) begin
    irqarray19_eventsourceflex306_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[2]) begin
        if (irqarray19_rising[2]) begin
            irqarray19_eventsourceflex306_trigger_filtered <= (irqarray19_interrupts[2] & (~irqarray19_eventsourceflex306_trigger_d));
        end else begin
            irqarray19_eventsourceflex306_trigger_filtered <= ((~irqarray19_interrupts[2]) & irqarray19_eventsourceflex306_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex306_trigger_filtered <= irqarray19_interrupts[2];
    end
end
assign irqarray19_eventsourceflex306_status = (irqarray19_interrupts[2] | irqarray19_trigger[2]);
always @(*) begin
    irqarray19_eventsourceflex307_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[3]) begin
        if (irqarray19_rising[3]) begin
            irqarray19_eventsourceflex307_trigger_filtered <= (irqarray19_interrupts[3] & (~irqarray19_eventsourceflex307_trigger_d));
        end else begin
            irqarray19_eventsourceflex307_trigger_filtered <= ((~irqarray19_interrupts[3]) & irqarray19_eventsourceflex307_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex307_trigger_filtered <= irqarray19_interrupts[3];
    end
end
assign irqarray19_eventsourceflex307_status = (irqarray19_interrupts[3] | irqarray19_trigger[3]);
always @(*) begin
    irqarray19_eventsourceflex308_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[4]) begin
        if (irqarray19_rising[4]) begin
            irqarray19_eventsourceflex308_trigger_filtered <= (irqarray19_interrupts[4] & (~irqarray19_eventsourceflex308_trigger_d));
        end else begin
            irqarray19_eventsourceflex308_trigger_filtered <= ((~irqarray19_interrupts[4]) & irqarray19_eventsourceflex308_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex308_trigger_filtered <= irqarray19_interrupts[4];
    end
end
assign irqarray19_eventsourceflex308_status = (irqarray19_interrupts[4] | irqarray19_trigger[4]);
always @(*) begin
    irqarray19_eventsourceflex309_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[5]) begin
        if (irqarray19_rising[5]) begin
            irqarray19_eventsourceflex309_trigger_filtered <= (irqarray19_interrupts[5] & (~irqarray19_eventsourceflex309_trigger_d));
        end else begin
            irqarray19_eventsourceflex309_trigger_filtered <= ((~irqarray19_interrupts[5]) & irqarray19_eventsourceflex309_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex309_trigger_filtered <= irqarray19_interrupts[5];
    end
end
assign irqarray19_eventsourceflex309_status = (irqarray19_interrupts[5] | irqarray19_trigger[5]);
always @(*) begin
    irqarray19_eventsourceflex310_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[6]) begin
        if (irqarray19_rising[6]) begin
            irqarray19_eventsourceflex310_trigger_filtered <= (irqarray19_interrupts[6] & (~irqarray19_eventsourceflex310_trigger_d));
        end else begin
            irqarray19_eventsourceflex310_trigger_filtered <= ((~irqarray19_interrupts[6]) & irqarray19_eventsourceflex310_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex310_trigger_filtered <= irqarray19_interrupts[6];
    end
end
assign irqarray19_eventsourceflex310_status = (irqarray19_interrupts[6] | irqarray19_trigger[6]);
always @(*) begin
    irqarray19_eventsourceflex311_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[7]) begin
        if (irqarray19_rising[7]) begin
            irqarray19_eventsourceflex311_trigger_filtered <= (irqarray19_interrupts[7] & (~irqarray19_eventsourceflex311_trigger_d));
        end else begin
            irqarray19_eventsourceflex311_trigger_filtered <= ((~irqarray19_interrupts[7]) & irqarray19_eventsourceflex311_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex311_trigger_filtered <= irqarray19_interrupts[7];
    end
end
assign irqarray19_eventsourceflex311_status = (irqarray19_interrupts[7] | irqarray19_trigger[7]);
always @(*) begin
    irqarray19_eventsourceflex312_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[8]) begin
        if (irqarray19_rising[8]) begin
            irqarray19_eventsourceflex312_trigger_filtered <= (irqarray19_interrupts[8] & (~irqarray19_eventsourceflex312_trigger_d));
        end else begin
            irqarray19_eventsourceflex312_trigger_filtered <= ((~irqarray19_interrupts[8]) & irqarray19_eventsourceflex312_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex312_trigger_filtered <= irqarray19_interrupts[8];
    end
end
assign irqarray19_eventsourceflex312_status = (irqarray19_interrupts[8] | irqarray19_trigger[8]);
always @(*) begin
    irqarray19_eventsourceflex313_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[9]) begin
        if (irqarray19_rising[9]) begin
            irqarray19_eventsourceflex313_trigger_filtered <= (irqarray19_interrupts[9] & (~irqarray19_eventsourceflex313_trigger_d));
        end else begin
            irqarray19_eventsourceflex313_trigger_filtered <= ((~irqarray19_interrupts[9]) & irqarray19_eventsourceflex313_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex313_trigger_filtered <= irqarray19_interrupts[9];
    end
end
assign irqarray19_eventsourceflex313_status = (irqarray19_interrupts[9] | irqarray19_trigger[9]);
always @(*) begin
    irqarray19_eventsourceflex314_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[10]) begin
        if (irqarray19_rising[10]) begin
            irqarray19_eventsourceflex314_trigger_filtered <= (irqarray19_interrupts[10] & (~irqarray19_eventsourceflex314_trigger_d));
        end else begin
            irqarray19_eventsourceflex314_trigger_filtered <= ((~irqarray19_interrupts[10]) & irqarray19_eventsourceflex314_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex314_trigger_filtered <= irqarray19_interrupts[10];
    end
end
assign irqarray19_eventsourceflex314_status = (irqarray19_interrupts[10] | irqarray19_trigger[10]);
always @(*) begin
    irqarray19_eventsourceflex315_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[11]) begin
        if (irqarray19_rising[11]) begin
            irqarray19_eventsourceflex315_trigger_filtered <= (irqarray19_interrupts[11] & (~irqarray19_eventsourceflex315_trigger_d));
        end else begin
            irqarray19_eventsourceflex315_trigger_filtered <= ((~irqarray19_interrupts[11]) & irqarray19_eventsourceflex315_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex315_trigger_filtered <= irqarray19_interrupts[11];
    end
end
assign irqarray19_eventsourceflex315_status = (irqarray19_interrupts[11] | irqarray19_trigger[11]);
always @(*) begin
    irqarray19_eventsourceflex316_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[12]) begin
        if (irqarray19_rising[12]) begin
            irqarray19_eventsourceflex316_trigger_filtered <= (irqarray19_interrupts[12] & (~irqarray19_eventsourceflex316_trigger_d));
        end else begin
            irqarray19_eventsourceflex316_trigger_filtered <= ((~irqarray19_interrupts[12]) & irqarray19_eventsourceflex316_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex316_trigger_filtered <= irqarray19_interrupts[12];
    end
end
assign irqarray19_eventsourceflex316_status = (irqarray19_interrupts[12] | irqarray19_trigger[12]);
always @(*) begin
    irqarray19_eventsourceflex317_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[13]) begin
        if (irqarray19_rising[13]) begin
            irqarray19_eventsourceflex317_trigger_filtered <= (irqarray19_interrupts[13] & (~irqarray19_eventsourceflex317_trigger_d));
        end else begin
            irqarray19_eventsourceflex317_trigger_filtered <= ((~irqarray19_interrupts[13]) & irqarray19_eventsourceflex317_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex317_trigger_filtered <= irqarray19_interrupts[13];
    end
end
assign irqarray19_eventsourceflex317_status = (irqarray19_interrupts[13] | irqarray19_trigger[13]);
always @(*) begin
    irqarray19_eventsourceflex318_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[14]) begin
        if (irqarray19_rising[14]) begin
            irqarray19_eventsourceflex318_trigger_filtered <= (irqarray19_interrupts[14] & (~irqarray19_eventsourceflex318_trigger_d));
        end else begin
            irqarray19_eventsourceflex318_trigger_filtered <= ((~irqarray19_interrupts[14]) & irqarray19_eventsourceflex318_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex318_trigger_filtered <= irqarray19_interrupts[14];
    end
end
assign irqarray19_eventsourceflex318_status = (irqarray19_interrupts[14] | irqarray19_trigger[14]);
always @(*) begin
    irqarray19_eventsourceflex319_trigger_filtered <= 1'd0;
    if (irqarray19_use_edge[15]) begin
        if (irqarray19_rising[15]) begin
            irqarray19_eventsourceflex319_trigger_filtered <= (irqarray19_interrupts[15] & (~irqarray19_eventsourceflex319_trigger_d));
        end else begin
            irqarray19_eventsourceflex319_trigger_filtered <= ((~irqarray19_interrupts[15]) & irqarray19_eventsourceflex319_trigger_d);
        end
    end else begin
        irqarray19_eventsourceflex319_trigger_filtered <= irqarray19_interrupts[15];
    end
end
assign irqarray19_eventsourceflex319_status = (irqarray19_interrupts[15] | irqarray19_trigger[15]);
assign ticktimer_load_xfer_i = ticktimer_load;
assign ticktimer_timer_sync_i = ticktimer_timer0;
assign ticktimer_timer1 = ticktimer_timer_sync_o;
assign ticktimer_resume_sync_i = ticktimer_resume_time;
assign ticktimer_time_status = ticktimer_timer_sync_o;
assign ticktimer_reset_xfer_i = ticktimer_reset;
assign ticktimer_alarm_trigger0 = ticktimer_alarm_trigger1;
assign ticktimer_ping_i = ticktimer_msleep_target_re;
assign ticktimer_pong_i = ticktimer_ping_o;
always @(*) begin
    ticktimer_alarm_trigger1 <= 1'd0;
    if (ticktimer_lockout_alarm) begin
        ticktimer_alarm_trigger1 <= 1'd0;
    end else begin
        ticktimer_alarm_trigger1 <= (ticktimer_msleep_target_storage <= ticktimer_timer_sync_o);
    end
end
assign ticktimer_target_xfer_i = ticktimer_msleep_target_storage;
assign ticktimer_alarm_always_on = ticktimer_alarm3;
assign ticktimer_clkspertick = ticktimer_clocks_per_tick_storage;
assign ticktimer_load_xfer_ps_i = (ticktimer_load_xfer_i & (~ticktimer_load_xfer_blind));
assign ticktimer_load_xfer_ps_ack_i = ticktimer_load_xfer_ps_o;
assign ticktimer_load_xfer_o = ticktimer_load_xfer_ps_o;
assign ticktimer_load_xfer_ps_o = (ticktimer_load_xfer_ps_toggle_o ^ ticktimer_load_xfer_ps_toggle_o_r);
assign ticktimer_load_xfer_ps_ack_o = (ticktimer_load_xfer_ps_ack_toggle_o ^ ticktimer_load_xfer_ps_ack_toggle_o_r);
assign ticktimer_timer_sync_wait = (~ticktimer_timer_sync_ping_i);
assign ticktimer_timer_sync_ping_i = ((ticktimer_timer_sync_starter | ticktimer_timer_sync_pong_o) | ticktimer_timer_sync_done);
assign ticktimer_timer_sync_pong_i = ticktimer_timer_sync_ping_o1;
assign ticktimer_timer_sync_ping_o0 = (ticktimer_timer_sync_ping_toggle_o ^ ticktimer_timer_sync_ping_toggle_o_r);
assign ticktimer_timer_sync_pong_o = (ticktimer_timer_sync_pong_toggle_o ^ ticktimer_timer_sync_pong_toggle_o_r);
assign ticktimer_timer_sync_done = (ticktimer_timer_sync_count == 1'd0);
assign ticktimer_resume_sync_wait = (~ticktimer_resume_sync_ping_i);
assign ticktimer_resume_sync_ping_i = ((ticktimer_resume_sync_starter | ticktimer_resume_sync_pong_o) | ticktimer_resume_sync_done);
assign ticktimer_resume_sync_pong_i = ticktimer_resume_sync_ping_o1;
assign ticktimer_resume_sync_ping_o0 = (ticktimer_resume_sync_ping_toggle_o ^ ticktimer_resume_sync_ping_toggle_o_r);
assign ticktimer_resume_sync_pong_o = (ticktimer_resume_sync_pong_toggle_o ^ ticktimer_resume_sync_pong_toggle_o_r);
assign ticktimer_resume_sync_done = (ticktimer_resume_sync_count == 1'd0);
assign ticktimer_reset_xfer_ps_i = (ticktimer_reset_xfer_i & (~ticktimer_reset_xfer_blind));
assign ticktimer_reset_xfer_ps_ack_i = ticktimer_reset_xfer_ps_o;
assign ticktimer_reset_xfer_o = ticktimer_reset_xfer_ps_o;
assign ticktimer_reset_xfer_ps_o = (ticktimer_reset_xfer_ps_toggle_o ^ ticktimer_reset_xfer_ps_toggle_o_r);
assign ticktimer_reset_xfer_ps_ack_o = (ticktimer_reset_xfer_ps_ack_toggle_o ^ ticktimer_reset_xfer_ps_ack_toggle_o_r);
assign ticktimer_alarm0 = ticktimer_alarm_status;
assign ticktimer_alarm1 = ticktimer_alarm_pending;
always @(*) begin
    ticktimer_alarm_clear <= 1'd0;
    if ((ticktimer_pending_re & ticktimer_pending_r)) begin
        ticktimer_alarm_clear <= 1'd1;
    end
end
assign ticktimer_irq = (ticktimer_pending_status & ticktimer_enable_storage);
assign ticktimer_alarm_status = ticktimer_alarm_trigger0;
assign ticktimer_alarm_pending = ticktimer_alarm_trigger0;
assign ticktimer_ping_ps_i = (ticktimer_ping_i & (~ticktimer_ping_blind));
assign ticktimer_ping_ps_ack_i = ticktimer_ping_ps_o;
assign ticktimer_ping_o = ticktimer_ping_ps_o;
assign ticktimer_ping_ps_o = (ticktimer_ping_ps_toggle_o ^ ticktimer_ping_ps_toggle_o_r);
assign ticktimer_ping_ps_ack_o = (ticktimer_ping_ps_ack_toggle_o ^ ticktimer_ping_ps_ack_toggle_o_r);
assign ticktimer_pong_ps_i = (ticktimer_pong_i & (~ticktimer_pong_blind));
assign ticktimer_pong_ps_ack_i = ticktimer_pong_ps_o;
assign ticktimer_pong_o = ticktimer_pong_ps_o;
assign ticktimer_pong_ps_o = (ticktimer_pong_ps_toggle_o ^ ticktimer_pong_ps_toggle_o_r);
assign ticktimer_pong_ps_ack_o = (ticktimer_pong_ps_ack_toggle_o ^ ticktimer_pong_ps_ack_toggle_o_r);
assign ticktimer_target_xfer_wait = (~ticktimer_target_xfer_ping_i);
assign ticktimer_target_xfer_ping_i = ((ticktimer_target_xfer_starter | ticktimer_target_xfer_pong_o) | ticktimer_target_xfer_done);
assign ticktimer_target_xfer_pong_i = ticktimer_target_xfer_ping_o1;
assign ticktimer_target_xfer_ping_o0 = (ticktimer_target_xfer_ping_toggle_o ^ ticktimer_target_xfer_ping_toggle_o_r);
assign ticktimer_target_xfer_pong_o = (ticktimer_target_xfer_pong_toggle_o ^ ticktimer_target_xfer_pong_toggle_o_r);
assign ticktimer_target_xfer_done = (ticktimer_target_xfer_count == 1'd0);
assign d11ctime_beat = d11ctime_heartbeat;
assign susres_resume1 = susres_resume0;
assign susres_soft_int_trigger = (susres_interrupt | susres_kernel_resume_interrupt);
assign susres_soft_int0 = susres_soft_int_status;
assign susres_soft_int1 = susres_soft_int_pending;
always @(*) begin
    susres_soft_int_clear <= 1'd0;
    if ((susres_pending_re & susres_pending_r)) begin
        susres_soft_int_clear <= 1'd1;
    end
end
assign susres_irq = (susres_pending_status & susres_enable_storage);
assign susres_soft_int_status = susres_soft_int_trigger;
assign mailbox_error_trigger = (mailbox_tx_err | mailbox_rx_err);
assign mailbox_w_fifo_reset_sys = ((~mailbox_reset_n) | mailbox_abort);
assign mailbox_tx_words = mailbox_syncfifobufferedmacro0_level;
assign mailbox_tx_err = mailbox_w_over_bit;
always @(*) begin
    mailbox_w_over_flag <= 1'd0;
    mailbox_syncfifobufferedmacro0_fifo_we <= 1'd0;
    if ((mailbox_wdata_re & (~mailbox_syncfifobufferedmacro0_fifo_writable))) begin
        mailbox_w_over_flag <= 1'd1;
    end else begin
        if ((~mailbox_abort_in_progress1)) begin
            mailbox_syncfifobufferedmacro0_fifo_we <= mailbox_wdata_re;
        end
    end
end
assign mailbox_w_over_clear = mailbox_status_we1;
assign mailbox_syncfifobufferedmacro0_fifo_din = mailbox_wdata_storage;
assign mailbox_w_dat = mailbox_syncfifobufferedmacro0_fifo_dout;
assign mailbox_w_valid = mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_readable;
assign mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_re = mailbox_w_ready;
assign mailbox_w_done = mailbox_done;
assign mailbox_syncfifobufferedmacro0_cmbist = mailbox_cmbist;
assign mailbox_syncfifobufferedmacro0_cmatpg = mailbox_cmatpg;
assign mailbox_syncfifobufferedmacro0_vexsramtrm = mailbox_vexsramtrm;
assign mailbox_r_fifo_reset_sys = ((~mailbox_reset_n) | mailbox_abort);
assign mailbox_rx_words = mailbox_syncfifobufferedmacro1_level;
assign mailbox_rx_err = mailbox_r_over_bit;
always @(*) begin
    mailbox_r_over_flag <= 1'd0;
    mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_re <= 1'd0;
    if ((mailbox_rdata_we & (~mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_readable))) begin
        mailbox_r_over_flag <= 1'd1;
    end else begin
        mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_re <= mailbox_rdata_we;
    end
end
assign mailbox_r_over_clear = mailbox_status_we1;
assign mailbox_syncfifobufferedmacro1_fifo_din = mailbox_r_dat;
assign mailbox_rdata_status = mailbox_syncfifobufferedmacro1_fifo_dout;
assign mailbox_r_ready = (mailbox_syncfifobufferedmacro1_fifo_writable & mailbox_r_valid);
assign mailbox_syncfifobufferedmacro1_fifo_we = ((mailbox_r_valid & mailbox_syncfifobufferedmacro1_fifo_writable) & (~mailbox_abort_in_progress1));
assign mailbox_available_trigger = mailbox_r_done;
assign mailbox_syncfifobufferedmacro1_cmbist = mailbox_cmbist;
assign mailbox_syncfifobufferedmacro1_cmatpg = mailbox_cmatpg;
assign mailbox_syncfifobufferedmacro1_vexsramtrm = mailbox_vexsramtrm;
assign mailbox_abort_in_progress0 = mailbox_abort_in_progress1;
assign mailbox_abort_ack0 = mailbox_abort_ack1;
assign mailbox_available0 = mailbox_available_status;
assign mailbox_available1 = mailbox_available_pending;
always @(*) begin
    mailbox_available_clear <= 1'd0;
    if ((mailbox_pending_re & mailbox_pending_r[0])) begin
        mailbox_available_clear <= 1'd1;
    end
end
assign mailbox_abort_init0 = mailbox_abort_init_status;
assign mailbox_abort_init1 = mailbox_abort_init_pending;
always @(*) begin
    mailbox_abort_init_clear <= 1'd0;
    if ((mailbox_pending_re & mailbox_pending_r[1])) begin
        mailbox_abort_init_clear <= 1'd1;
    end
end
assign mailbox_abort_done0 = mailbox_abort_done_status;
assign mailbox_abort_done1 = mailbox_abort_done_pending;
always @(*) begin
    mailbox_abort_done_clear <= 1'd0;
    if ((mailbox_pending_re & mailbox_pending_r[2])) begin
        mailbox_abort_done_clear <= 1'd1;
    end
end
assign mailbox_error0 = mailbox_error_status;
assign mailbox_error1 = mailbox_error_pending;
always @(*) begin
    mailbox_error_clear <= 1'd0;
    if ((mailbox_pending_re & mailbox_pending_r[3])) begin
        mailbox_error_clear <= 1'd1;
    end
end
assign mailbox_irq = ((((mailbox_pending_status[0] & mailbox_enable_storage[0]) | (mailbox_pending_status[1] & mailbox_enable_storage[1])) | (mailbox_pending_status[2] & mailbox_enable_storage[2])) | (mailbox_pending_status[3] & mailbox_enable_storage[3]));
assign mailbox_available_status = 1'd0;
assign mailbox_abort_init_status = mailbox_abort_init_trigger;
assign mailbox_abort_done_status = mailbox_abort_done_trigger;
assign mailbox_error_status = mailbox_error_trigger;
assign mailbox_syncfifobufferedmacro0_fifo_cmbist = mailbox_syncfifobufferedmacro0_cmbist;
assign mailbox_syncfifobufferedmacro0_fifo_cmatpg = mailbox_syncfifobufferedmacro0_cmatpg;
assign mailbox_syncfifobufferedmacro0_fifo_vexsramtrm = mailbox_syncfifobufferedmacro0_vexsramtrm;
assign mailbox_syncfifobufferedmacro0_fifo_re = (mailbox_syncfifobufferedmacro0_fifo_readable & ((~mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_readable) | mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_re));
assign mailbox_syncfifobufferedmacro0_level = (mailbox_syncfifobufferedmacro0_fifo_level + mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_readable);
always @(*) begin
    mailbox_syncfifobufferedmacro0_fifo_wrport_adr <= 10'd0;
    if (1'd0) begin
        mailbox_syncfifobufferedmacro0_fifo_wrport_adr <= (mailbox_syncfifobufferedmacro0_fifo_produce - 1'd1);
    end else begin
        mailbox_syncfifobufferedmacro0_fifo_wrport_adr <= mailbox_syncfifobufferedmacro0_fifo_produce;
    end
end
assign mailbox_syncfifobufferedmacro0_fifo_wrport_dat_w = mailbox_syncfifobufferedmacro0_fifo_din;
assign mailbox_syncfifobufferedmacro0_fifo_wrport_we = (mailbox_syncfifobufferedmacro0_fifo_we & (mailbox_syncfifobufferedmacro0_fifo_writable | 1'd0));
assign mailbox_syncfifobufferedmacro0_fifo_do_read = (mailbox_syncfifobufferedmacro0_fifo_readable & mailbox_syncfifobufferedmacro0_fifo_re);
assign mailbox_syncfifobufferedmacro0_fifo_rdport_adr = mailbox_syncfifobufferedmacro0_fifo_consume;
assign mailbox_syncfifobufferedmacro0_fifo_dout = mailbox_syncfifobufferedmacro0_fifo_rdport_dat_r;
assign mailbox_syncfifobufferedmacro0_fifo_rdport_re = mailbox_syncfifobufferedmacro0_fifo_do_read;
assign mailbox_syncfifobufferedmacro0_fifo_writable = (mailbox_syncfifobufferedmacro0_fifo_level != 11'd1024);
assign mailbox_syncfifobufferedmacro0_fifo_readable = (mailbox_syncfifobufferedmacro0_fifo_level != 1'd0);
assign mailbox_syncfifobufferedmacro1_fifo_cmbist = mailbox_syncfifobufferedmacro1_cmbist;
assign mailbox_syncfifobufferedmacro1_fifo_cmatpg = mailbox_syncfifobufferedmacro1_cmatpg;
assign mailbox_syncfifobufferedmacro1_fifo_vexsramtrm = mailbox_syncfifobufferedmacro1_vexsramtrm;
assign mailbox_syncfifobufferedmacro1_fifo_re = (mailbox_syncfifobufferedmacro1_fifo_readable & ((~mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_readable) | mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_re));
assign mailbox_syncfifobufferedmacro1_level = (mailbox_syncfifobufferedmacro1_fifo_level + mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_readable);
always @(*) begin
    mailbox_syncfifobufferedmacro1_fifo_wrport_adr <= 10'd0;
    if (1'd0) begin
        mailbox_syncfifobufferedmacro1_fifo_wrport_adr <= (mailbox_syncfifobufferedmacro1_fifo_produce - 1'd1);
    end else begin
        mailbox_syncfifobufferedmacro1_fifo_wrport_adr <= mailbox_syncfifobufferedmacro1_fifo_produce;
    end
end
assign mailbox_syncfifobufferedmacro1_fifo_wrport_dat_w = mailbox_syncfifobufferedmacro1_fifo_din;
assign mailbox_syncfifobufferedmacro1_fifo_wrport_we = (mailbox_syncfifobufferedmacro1_fifo_we & (mailbox_syncfifobufferedmacro1_fifo_writable | 1'd0));
assign mailbox_syncfifobufferedmacro1_fifo_do_read = (mailbox_syncfifobufferedmacro1_fifo_readable & mailbox_syncfifobufferedmacro1_fifo_re);
assign mailbox_syncfifobufferedmacro1_fifo_rdport_adr = mailbox_syncfifobufferedmacro1_fifo_consume;
assign mailbox_syncfifobufferedmacro1_fifo_dout = mailbox_syncfifobufferedmacro1_fifo_rdport_dat_r;
assign mailbox_syncfifobufferedmacro1_fifo_rdport_re = mailbox_syncfifobufferedmacro1_fifo_do_read;
assign mailbox_syncfifobufferedmacro1_fifo_writable = (mailbox_syncfifobufferedmacro1_fifo_level != 11'd1024);
assign mailbox_syncfifobufferedmacro1_fifo_readable = (mailbox_syncfifobufferedmacro1_fifo_level != 1'd0);
always @(*) begin
    cramsoc_mailbox_next_state <= 2'd0;
    mailbox_abort_ack1_mailbox_next_value0 <= 1'd0;
    mailbox_abort_done_trigger <= 1'd0;
    mailbox_abort_ack1_mailbox_next_value_ce0 <= 1'd0;
    mailbox_abort_in_progress1_mailbox_next_value1 <= 1'd0;
    mailbox_abort_in_progress1_mailbox_next_value_ce1 <= 1'd0;
    mailbox_w_abort_mailbox_next_value2 <= 1'd0;
    mailbox_w_abort_mailbox_next_value_ce2 <= 1'd0;
    mailbox_abort_init_trigger <= 1'd0;
    cramsoc_mailbox_next_state <= cramsoc_mailbox_state;
    case (cramsoc_mailbox_state)
        1'd1: begin
            if (mailbox_r_abort) begin
                cramsoc_mailbox_next_state <= 1'd0;
                mailbox_abort_in_progress1_mailbox_next_value1 <= 1'd0;
                mailbox_abort_in_progress1_mailbox_next_value_ce1 <= 1'd1;
                mailbox_abort_done_trigger <= 1'd1;
                mailbox_w_abort_mailbox_next_value2 <= 1'd0;
                mailbox_w_abort_mailbox_next_value_ce2 <= 1'd1;
            end else begin
                mailbox_w_abort_mailbox_next_value2 <= 1'd1;
                mailbox_w_abort_mailbox_next_value_ce2 <= 1'd1;
            end
        end
        2'd2: begin
            if (mailbox_abort) begin
                cramsoc_mailbox_next_state <= 2'd3;
                mailbox_abort_in_progress1_mailbox_next_value1 <= 1'd0;
                mailbox_abort_in_progress1_mailbox_next_value_ce1 <= 1'd1;
                mailbox_abort_ack1_mailbox_next_value0 <= 1'd1;
                mailbox_abort_ack1_mailbox_next_value_ce0 <= 1'd1;
                mailbox_w_abort_mailbox_next_value2 <= 1'd1;
                mailbox_w_abort_mailbox_next_value_ce2 <= 1'd1;
            end
        end
        2'd3: begin
            cramsoc_mailbox_next_state <= 1'd0;
            mailbox_w_abort_mailbox_next_value2 <= 1'd0;
            mailbox_w_abort_mailbox_next_value_ce2 <= 1'd1;
        end
        default: begin
            if ((mailbox_abort & (~mailbox_r_abort))) begin
                cramsoc_mailbox_next_state <= 1'd1;
                mailbox_abort_ack1_mailbox_next_value0 <= 1'd0;
                mailbox_abort_ack1_mailbox_next_value_ce0 <= 1'd1;
                mailbox_abort_in_progress1_mailbox_next_value1 <= 1'd1;
                mailbox_abort_in_progress1_mailbox_next_value_ce1 <= 1'd1;
                mailbox_w_abort_mailbox_next_value2 <= 1'd1;
                mailbox_w_abort_mailbox_next_value_ce2 <= 1'd1;
            end else begin
                if ((mailbox_abort & mailbox_r_abort)) begin
                    cramsoc_mailbox_next_state <= 1'd0;
                    mailbox_abort_ack1_mailbox_next_value0 <= 1'd1;
                    mailbox_abort_ack1_mailbox_next_value_ce0 <= 1'd1;
                    mailbox_w_abort_mailbox_next_value2 <= 1'd1;
                    mailbox_w_abort_mailbox_next_value_ce2 <= 1'd1;
                end else begin
                    if (((~mailbox_abort) & mailbox_r_abort)) begin
                        cramsoc_mailbox_next_state <= 2'd2;
                        mailbox_abort_in_progress1_mailbox_next_value1 <= 1'd1;
                        mailbox_abort_in_progress1_mailbox_next_value_ce1 <= 1'd1;
                        mailbox_abort_init_trigger <= 1'd1;
                        mailbox_w_abort_mailbox_next_value2 <= 1'd0;
                        mailbox_w_abort_mailbox_next_value_ce2 <= 1'd1;
                    end else begin
                        mailbox_w_abort_mailbox_next_value2 <= 1'd0;
                        mailbox_w_abort_mailbox_next_value_ce2 <= 1'd1;
                    end
                end
            end
        end
    endcase
end
assign mb_client_error_trigger = (mb_client_tx_err | mb_client_rx_err);
assign mb_client_w_dat = mb_client_wdata_storage;
assign mb_client_w_valid = (mb_client_wdata_re | mb_client_w_pending);
assign mb_client_w_done = mb_client_done;
assign mb_client_tx_free = (~(mb_client_w_valid | mb_client_w_pending));
assign mb_client_rdata_status = mb_client_r_dat;
assign mb_client_r_ready = mb_client_rdata_we;
assign mb_client_available_trigger = mb_client_r_done;
assign mb_client_rx_avail = mb_client_r_valid;
assign mb_client_abort_in_progress0 = mb_client_abort_in_progress1;
assign mb_client_abort_ack0 = mb_client_abort_ack1;
assign mb_client_available0 = mb_client_available_status;
assign mb_client_available1 = mb_client_available_pending;
always @(*) begin
    mb_client_available_clear <= 1'd0;
    if ((mb_client_pending_re & mb_client_pending_r[0])) begin
        mb_client_available_clear <= 1'd1;
    end
end
assign mb_client_abort_init0 = mb_client_abort_init_status;
assign mb_client_abort_init1 = mb_client_abort_init_pending;
always @(*) begin
    mb_client_abort_init_clear <= 1'd0;
    if ((mb_client_pending_re & mb_client_pending_r[1])) begin
        mb_client_abort_init_clear <= 1'd1;
    end
end
assign mb_client_abort_done0 = mb_client_abort_done_status;
assign mb_client_abort_done1 = mb_client_abort_done_pending;
always @(*) begin
    mb_client_abort_done_clear <= 1'd0;
    if ((mb_client_pending_re & mb_client_pending_r[2])) begin
        mb_client_abort_done_clear <= 1'd1;
    end
end
assign mb_client_error0 = mb_client_error_status;
assign mb_client_error1 = mb_client_error_pending;
always @(*) begin
    mb_client_error_clear <= 1'd0;
    if ((mb_client_pending_re & mb_client_pending_r[3])) begin
        mb_client_error_clear <= 1'd1;
    end
end
assign mb_client_irq = ((((mb_client_pending_status[0] & mb_client_enable_storage[0]) | (mb_client_pending_status[1] & mb_client_enable_storage[1])) | (mb_client_pending_status[2] & mb_client_enable_storage[2])) | (mb_client_pending_status[3] & mb_client_enable_storage[3]));
assign mb_client_available_status = 1'd0;
assign mb_client_abort_init_status = mb_client_abort_init_trigger;
assign mb_client_abort_done_status = mb_client_abort_done_trigger;
assign mb_client_error_status = mb_client_error_trigger;
always @(*) begin
    cramsoc_mailboxclient_next_state <= 2'd0;
    mb_client_abort_done_trigger <= 1'd0;
    mb_client_abort_ack1_mailboxclient_next_value0 <= 1'd0;
    mb_client_abort_ack1_mailboxclient_next_value_ce0 <= 1'd0;
    mb_client_abort_in_progress1_mailboxclient_next_value1 <= 1'd0;
    mb_client_abort_in_progress1_mailboxclient_next_value_ce1 <= 1'd0;
    mb_client_w_abort_mailboxclient_next_value2 <= 1'd0;
    mb_client_abort_init_trigger <= 1'd0;
    mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd0;
    cramsoc_mailboxclient_next_state <= cramsoc_mailboxclient_state;
    case (cramsoc_mailboxclient_state)
        1'd1: begin
            if (mb_client_r_abort) begin
                cramsoc_mailboxclient_next_state <= 1'd0;
                mb_client_abort_in_progress1_mailboxclient_next_value1 <= 1'd0;
                mb_client_abort_in_progress1_mailboxclient_next_value_ce1 <= 1'd1;
                mb_client_abort_done_trigger <= 1'd1;
                mb_client_w_abort_mailboxclient_next_value2 <= 1'd0;
                mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd1;
            end else begin
                mb_client_w_abort_mailboxclient_next_value2 <= 1'd1;
                mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd1;
            end
        end
        2'd2: begin
            if (mb_client_abort) begin
                cramsoc_mailboxclient_next_state <= 2'd3;
                mb_client_abort_in_progress1_mailboxclient_next_value1 <= 1'd0;
                mb_client_abort_in_progress1_mailboxclient_next_value_ce1 <= 1'd1;
                mb_client_abort_ack1_mailboxclient_next_value0 <= 1'd1;
                mb_client_abort_ack1_mailboxclient_next_value_ce0 <= 1'd1;
                mb_client_w_abort_mailboxclient_next_value2 <= 1'd1;
                mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd1;
            end
        end
        2'd3: begin
            cramsoc_mailboxclient_next_state <= 1'd0;
            mb_client_w_abort_mailboxclient_next_value2 <= 1'd0;
            mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd1;
        end
        default: begin
            if ((mb_client_abort & (~mb_client_r_abort))) begin
                cramsoc_mailboxclient_next_state <= 1'd1;
                mb_client_abort_ack1_mailboxclient_next_value0 <= 1'd0;
                mb_client_abort_ack1_mailboxclient_next_value_ce0 <= 1'd1;
                mb_client_abort_in_progress1_mailboxclient_next_value1 <= 1'd1;
                mb_client_abort_in_progress1_mailboxclient_next_value_ce1 <= 1'd1;
                mb_client_w_abort_mailboxclient_next_value2 <= 1'd1;
                mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd1;
            end else begin
                if ((mb_client_abort & mb_client_r_abort)) begin
                    cramsoc_mailboxclient_next_state <= 1'd0;
                    mb_client_abort_ack1_mailboxclient_next_value0 <= 1'd1;
                    mb_client_abort_ack1_mailboxclient_next_value_ce0 <= 1'd1;
                    mb_client_w_abort_mailboxclient_next_value2 <= 1'd1;
                    mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd1;
                end else begin
                    if (((~mb_client_abort) & mb_client_r_abort)) begin
                        cramsoc_mailboxclient_next_state <= 2'd2;
                        mb_client_abort_in_progress1_mailboxclient_next_value1 <= 1'd1;
                        mb_client_abort_in_progress1_mailboxclient_next_value_ce1 <= 1'd1;
                        mb_client_abort_init_trigger <= 1'd1;
                        mb_client_w_abort_mailboxclient_next_value2 <= 1'd0;
                        mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd1;
                    end else begin
                        mb_client_w_abort_mailboxclient_next_value2 <= 1'd0;
                        mb_client_w_abort_mailboxclient_next_value_ce2 <= 1'd1;
                    end
                end
            end
        end
    endcase
end
assign csr_rtest_status = (csr_wtest_storage + 29'd268435456);
assign cramsoc_dat_w = cramsoc_w_payload_data;
assign cramsoc_we = ((cramsoc_w_valid & cramsoc_w_ready) & (cramsoc_w_payload_strb != 1'd0));
assign cramsoc_re = cramsoc_r_ready;
always @(*) begin
    cramsoc_do_read <= 1'd0;
    cramsoc_do_write <= 1'd0;
    if ((cramsoc_aw_valid & cramsoc_ar_valid)) begin
        cramsoc_do_write <= cramsoc_last_was_read;
        cramsoc_do_read <= (~cramsoc_last_was_read);
    end else begin
        cramsoc_do_write <= cramsoc_aw_valid;
        cramsoc_do_read <= cramsoc_ar_valid;
    end
end
assign cramsoc_r_valid = cramsoc_nocomb_axl_r_valid;
assign cramsoc_aw_ready = cramsoc_nocomb_axl_aw_ready;
assign cramsoc_w_ready = cramsoc_nocomb_axl_w_ready;
assign cramsoc_ar_ready = cramsoc_nocomb_axl_ar_ready;
assign cramsoc_b_valid = cramsoc_nocomb_axl_b_valid;
always @(*) begin
    cramsoc_axilite2csr_next_state <= 2'd0;
    cramsoc_adr <= 16'd0;
    cramsoc_r_payload_data <= 32'd0;
    cramsoc_r_payload_resp <= 2'd0;
    cramsoc_last_was_read_axilite2csr_next_value <= 1'd0;
    cramsoc_last_was_read_axilite2csr_next_value_ce <= 1'd0;
    cramsoc_b_payload_resp <= 2'd0;
    cramsoc_nocomb_axl_r_valid <= 1'd0;
    cramsoc_nocomb_axl_w_ready <= 1'd0;
    cramsoc_nocomb_axl_aw_ready <= 1'd0;
    cramsoc_nocomb_axl_ar_ready <= 1'd0;
    cramsoc_nocomb_axl_b_valid <= 1'd0;
    cramsoc_axilite2csr_next_state <= cramsoc_axilite2csr_state;
    case (cramsoc_axilite2csr_state)
        1'd1: begin
            cramsoc_last_was_read_axilite2csr_next_value <= 1'd1;
            cramsoc_last_was_read_axilite2csr_next_value_ce <= 1'd1;
            cramsoc_adr <= cramsoc_ar_payload_addr[31:2];
            cramsoc_r_payload_data <= cramsoc_dat_r;
            cramsoc_r_payload_resp <= 1'd0;
            cramsoc_nocomb_axl_r_valid <= 1'd1;
            if (cramsoc_r_ready) begin
                cramsoc_axilite2csr_next_state <= 1'd0;
            end
        end
        2'd2: begin
            cramsoc_last_was_read_axilite2csr_next_value <= 1'd0;
            cramsoc_last_was_read_axilite2csr_next_value_ce <= 1'd1;
            cramsoc_nocomb_axl_b_valid <= 1'd1;
            cramsoc_b_payload_resp <= 1'd0;
            if (cramsoc_b_ready) begin
                cramsoc_axilite2csr_next_state <= 1'd0;
            end
        end
        default: begin
            if (cramsoc_do_write) begin
                cramsoc_adr <= cramsoc_aw_payload_addr[31:2];
                if (cramsoc_w_valid) begin
                    cramsoc_nocomb_axl_aw_ready <= 1'd1;
                    cramsoc_nocomb_axl_w_ready <= 1'd1;
                    cramsoc_axilite2csr_next_state <= 2'd2;
                end
            end else begin
                if (cramsoc_do_read) begin
                    cramsoc_nocomb_axl_ar_ready <= 1'd1;
                    cramsoc_adr <= cramsoc_ar_payload_addr[31:2];
                    cramsoc_axilite2csr_next_state <= 1'd1;
                end
            end
        end
    endcase
end
assign csrbank0_sel = (interface0_bank_bus_adr[15:10] == 2'd2);
assign csrbank0_re = interface0_bank_bus_re;
assign csrbank0_control0_r = interface0_bank_bus_dat_w[1:0];
always @(*) begin
    csrbank0_control0_re <= 1'd0;
    csrbank0_control0_we <= 1'd0;
    if ((csrbank0_sel & (interface0_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank0_control0_re <= interface0_bank_bus_we;
        csrbank0_control0_we <= csrbank0_re;
    end
end
assign csrbank0_status_r = interface0_bank_bus_dat_w[8:0];
always @(*) begin
    csrbank0_status_we <= 1'd0;
    csrbank0_status_re <= 1'd0;
    if ((csrbank0_sel & (interface0_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank0_status_re <= interface0_bank_bus_we;
        csrbank0_status_we <= csrbank0_re;
    end
end
assign csrbank0_map_lo0_r = interface0_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank0_map_lo0_we <= 1'd0;
    csrbank0_map_lo0_re <= 1'd0;
    if ((csrbank0_sel & (interface0_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank0_map_lo0_re <= interface0_bank_bus_we;
        csrbank0_map_lo0_we <= csrbank0_re;
    end
end
assign csrbank0_map_hi0_r = interface0_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank0_map_hi0_re <= 1'd0;
    csrbank0_map_hi0_we <= 1'd0;
    if ((csrbank0_sel & (interface0_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank0_map_hi0_re <= interface0_bank_bus_we;
        csrbank0_map_hi0_we <= csrbank0_re;
    end
end
assign csrbank0_uservalue0_r = interface0_bank_bus_dat_w[17:0];
always @(*) begin
    csrbank0_uservalue0_we <= 1'd0;
    csrbank0_uservalue0_re <= 1'd0;
    if ((csrbank0_sel & (interface0_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank0_uservalue0_re <= interface0_bank_bus_we;
        csrbank0_uservalue0_we <= csrbank0_re;
    end
end
assign csrbank0_protect0_r = interface0_bank_bus_dat_w[0];
always @(*) begin
    csrbank0_protect0_we <= 1'd0;
    csrbank0_protect0_re <= 1'd0;
    if ((csrbank0_sel & (interface0_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank0_protect0_re <= interface0_bank_bus_we;
        csrbank0_protect0_we <= csrbank0_re;
    end
end
assign coreuser_enable0 = coreuser_control_storage[0];
assign coreuser_invert_priv0 = coreuser_control_storage[1];
assign csrbank0_control0_w = coreuser_control_storage[1:0];
always @(*) begin
    coreuser_status_status <= 9'd0;
    coreuser_status_status[7:0] <= coreuser_coreuser;
    coreuser_status_status[8] <= coreuser_mm;
end
assign csrbank0_status_w = coreuser_status_status[8:0];
assign coreuser_status_we = csrbank0_status_we;
assign coreuser_lut00 = coreuser_map_lo_storage[7:0];
assign coreuser_lut10 = coreuser_map_lo_storage[15:8];
assign coreuser_lut20 = coreuser_map_lo_storage[23:16];
assign coreuser_lut30 = coreuser_map_lo_storage[31:24];
assign csrbank0_map_lo0_w = coreuser_map_lo_storage[31:0];
assign coreuser_lut40 = coreuser_map_hi_storage[7:0];
assign coreuser_lut50 = coreuser_map_hi_storage[15:8];
assign coreuser_lut60 = coreuser_map_hi_storage[23:16];
assign coreuser_lut70 = coreuser_map_hi_storage[31:24];
assign csrbank0_map_hi0_w = coreuser_map_hi_storage[31:0];
assign coreuser_user00 = coreuser_uservalue_storage[1:0];
assign coreuser_user10 = coreuser_uservalue_storage[3:2];
assign coreuser_user20 = coreuser_uservalue_storage[5:4];
assign coreuser_user30 = coreuser_uservalue_storage[7:6];
assign coreuser_user40 = coreuser_uservalue_storage[9:8];
assign coreuser_user50 = coreuser_uservalue_storage[11:10];
assign coreuser_user60 = coreuser_uservalue_storage[13:12];
assign coreuser_user70 = coreuser_uservalue_storage[15:14];
assign coreuser_default = coreuser_uservalue_storage[17:16];
assign csrbank0_uservalue0_w = coreuser_uservalue_storage[17:0];
assign csrbank0_protect0_w = coreuser_protect_storage;
assign csrbank1_sel = (interface1_bank_bus_adr[15:10] == 2'd3);
assign csrbank1_re = interface1_bank_bus_re;
assign csrbank1_wtest0_r = interface1_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank1_wtest0_re <= 1'd0;
    csrbank1_wtest0_we <= 1'd0;
    if ((csrbank1_sel & (interface1_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank1_wtest0_re <= interface1_bank_bus_we;
        csrbank1_wtest0_we <= csrbank1_re;
    end
end
assign csrbank1_rtest_r = interface1_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank1_rtest_we <= 1'd0;
    csrbank1_rtest_re <= 1'd0;
    if ((csrbank1_sel & (interface1_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank1_rtest_re <= interface1_bank_bus_we;
        csrbank1_rtest_we <= csrbank1_re;
    end
end
assign csrbank1_wtest0_w = csr_wtest_storage[31:0];
assign csrbank1_rtest_w = csr_rtest_status[31:0];
assign csr_rtest_we = csrbank1_rtest_we;
assign csrbank2_sel = (interface2_bank_bus_adr[15:10] == 1'd0);
assign csrbank2_re = interface2_bank_bus_re;
assign csrbank2_control0_r = interface2_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank2_control0_we <= 1'd0;
    csrbank2_control0_re <= 1'd0;
    if ((csrbank2_sel & (interface2_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank2_control0_re <= interface2_bank_bus_we;
        csrbank2_control0_we <= csrbank2_re;
    end
end
assign csrbank2_heartbeat_r = interface2_bank_bus_dat_w[0];
always @(*) begin
    csrbank2_heartbeat_re <= 1'd0;
    csrbank2_heartbeat_we <= 1'd0;
    if ((csrbank2_sel & (interface2_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank2_heartbeat_re <= interface2_bank_bus_we;
        csrbank2_heartbeat_we <= csrbank2_re;
    end
end
assign d11ctime_count = d11ctime_control_storage[31:0];
assign csrbank2_control0_w = d11ctime_control_storage[31:0];
assign d11ctime_heartbeat_status = d11ctime_beat;
assign csrbank2_heartbeat_w = d11ctime_heartbeat_status;
assign d11ctime_heartbeat_we = csrbank2_heartbeat_we;
assign csrbank3_sel = (interface3_bank_bus_adr[15:10] == 3'd4);
assign csrbank3_re = interface3_bank_bus_re;
assign csrbank3_ev_soft0_r = interface3_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank3_ev_soft0_re <= 1'd0;
    csrbank3_ev_soft0_we <= 1'd0;
    if ((csrbank3_sel & (interface3_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank3_ev_soft0_re <= interface3_bank_bus_we;
        csrbank3_ev_soft0_we <= csrbank3_re;
    end
end
assign csrbank3_ev_edge_triggered0_r = interface3_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank3_ev_edge_triggered0_we <= 1'd0;
    csrbank3_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank3_sel & (interface3_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank3_ev_edge_triggered0_re <= interface3_bank_bus_we;
        csrbank3_ev_edge_triggered0_we <= csrbank3_re;
    end
end
assign csrbank3_ev_polarity0_r = interface3_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank3_ev_polarity0_we <= 1'd0;
    csrbank3_ev_polarity0_re <= 1'd0;
    if ((csrbank3_sel & (interface3_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank3_ev_polarity0_re <= interface3_bank_bus_we;
        csrbank3_ev_polarity0_we <= csrbank3_re;
    end
end
assign csrbank3_ev_status_r = interface3_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank3_ev_status_re <= 1'd0;
    csrbank3_ev_status_we <= 1'd0;
    if ((csrbank3_sel & (interface3_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank3_ev_status_re <= interface3_bank_bus_we;
        csrbank3_ev_status_we <= csrbank3_re;
    end
end
assign csrbank3_ev_pending_r = interface3_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank3_ev_pending_we <= 1'd0;
    csrbank3_ev_pending_re <= 1'd0;
    if ((csrbank3_sel & (interface3_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank3_ev_pending_re <= interface3_bank_bus_we;
        csrbank3_ev_pending_we <= csrbank3_re;
    end
end
assign csrbank3_ev_enable0_r = interface3_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank3_ev_enable0_we <= 1'd0;
    csrbank3_ev_enable0_re <= 1'd0;
    if ((csrbank3_sel & (interface3_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank3_ev_enable0_re <= interface3_bank_bus_we;
        csrbank3_ev_enable0_we <= csrbank3_re;
    end
end
always @(*) begin
    irqarray0_trigger <= 16'd0;
    if (irqarray0_soft_re) begin
        irqarray0_trigger <= irqarray0_soft_storage[15:0];
    end
end
assign csrbank3_ev_soft0_w = irqarray0_soft_storage[15:0];
assign irqarray0_use_edge = irqarray0_edge_triggered_storage[15:0];
assign csrbank3_ev_edge_triggered0_w = irqarray0_edge_triggered_storage[15:0];
assign irqarray0_rising = irqarray0_polarity_storage[15:0];
assign csrbank3_ev_polarity0_w = irqarray0_polarity_storage[15:0];
always @(*) begin
    irqarray0_status_status <= 16'd0;
    irqarray0_status_status[0] <= irqarray0_mdmairq_dupe0;
    irqarray0_status_status[1] <= irqarray0_nc_b0s10;
    irqarray0_status_status[2] <= irqarray0_nc_b0s20;
    irqarray0_status_status[3] <= irqarray0_nc_b0s30;
    irqarray0_status_status[4] <= irqarray0_pioirq0_dupe0;
    irqarray0_status_status[5] <= irqarray0_pioirq1_dupe0;
    irqarray0_status_status[6] <= irqarray0_pioirq2_dupe0;
    irqarray0_status_status[7] <= irqarray0_pioirq3_dupe0;
    irqarray0_status_status[8] <= irqarray0_nc_b0s80;
    irqarray0_status_status[9] <= irqarray0_nc_b0s90;
    irqarray0_status_status[10] <= irqarray0_nc_b0s100;
    irqarray0_status_status[11] <= irqarray0_nc_b0s110;
    irqarray0_status_status[12] <= irqarray0_nc_b0s120;
    irqarray0_status_status[13] <= irqarray0_nc_b0s130;
    irqarray0_status_status[14] <= irqarray0_nc_b0s140;
    irqarray0_status_status[15] <= irqarray0_nc_b0s150;
end
assign csrbank3_ev_status_w = irqarray0_status_status[15:0];
assign irqarray0_status_we = csrbank3_ev_status_we;
always @(*) begin
    irqarray0_pending_status <= 16'd0;
    irqarray0_pending_status[0] <= irqarray0_mdmairq_dupe1;
    irqarray0_pending_status[1] <= irqarray0_nc_b0s11;
    irqarray0_pending_status[2] <= irqarray0_nc_b0s21;
    irqarray0_pending_status[3] <= irqarray0_nc_b0s31;
    irqarray0_pending_status[4] <= irqarray0_pioirq0_dupe1;
    irqarray0_pending_status[5] <= irqarray0_pioirq1_dupe1;
    irqarray0_pending_status[6] <= irqarray0_pioirq2_dupe1;
    irqarray0_pending_status[7] <= irqarray0_pioirq3_dupe1;
    irqarray0_pending_status[8] <= irqarray0_nc_b0s81;
    irqarray0_pending_status[9] <= irqarray0_nc_b0s91;
    irqarray0_pending_status[10] <= irqarray0_nc_b0s101;
    irqarray0_pending_status[11] <= irqarray0_nc_b0s111;
    irqarray0_pending_status[12] <= irqarray0_nc_b0s121;
    irqarray0_pending_status[13] <= irqarray0_nc_b0s131;
    irqarray0_pending_status[14] <= irqarray0_nc_b0s141;
    irqarray0_pending_status[15] <= irqarray0_nc_b0s151;
end
assign csrbank3_ev_pending_w = irqarray0_pending_status[15:0];
assign irqarray0_pending_we = csrbank3_ev_pending_we;
assign irqarray0_mdmairq_dupe2 = irqarray0_enable_storage[0];
assign irqarray0_nc_b0s12 = irqarray0_enable_storage[1];
assign irqarray0_nc_b0s22 = irqarray0_enable_storage[2];
assign irqarray0_nc_b0s32 = irqarray0_enable_storage[3];
assign irqarray0_pioirq0_dupe2 = irqarray0_enable_storage[4];
assign irqarray0_pioirq1_dupe2 = irqarray0_enable_storage[5];
assign irqarray0_pioirq2_dupe2 = irqarray0_enable_storage[6];
assign irqarray0_pioirq3_dupe2 = irqarray0_enable_storage[7];
assign irqarray0_nc_b0s82 = irqarray0_enable_storage[8];
assign irqarray0_nc_b0s92 = irqarray0_enable_storage[9];
assign irqarray0_nc_b0s102 = irqarray0_enable_storage[10];
assign irqarray0_nc_b0s112 = irqarray0_enable_storage[11];
assign irqarray0_nc_b0s122 = irqarray0_enable_storage[12];
assign irqarray0_nc_b0s132 = irqarray0_enable_storage[13];
assign irqarray0_nc_b0s142 = irqarray0_enable_storage[14];
assign irqarray0_nc_b0s152 = irqarray0_enable_storage[15];
assign csrbank3_ev_enable0_w = irqarray0_enable_storage[15:0];
assign csrbank4_sel = (interface4_bank_bus_adr[15:10] == 3'd5);
assign csrbank4_re = interface4_bank_bus_re;
assign csrbank4_ev_soft0_r = interface4_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank4_ev_soft0_re <= 1'd0;
    csrbank4_ev_soft0_we <= 1'd0;
    if ((csrbank4_sel & (interface4_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank4_ev_soft0_re <= interface4_bank_bus_we;
        csrbank4_ev_soft0_we <= csrbank4_re;
    end
end
assign csrbank4_ev_edge_triggered0_r = interface4_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank4_ev_edge_triggered0_we <= 1'd0;
    csrbank4_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank4_sel & (interface4_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank4_ev_edge_triggered0_re <= interface4_bank_bus_we;
        csrbank4_ev_edge_triggered0_we <= csrbank4_re;
    end
end
assign csrbank4_ev_polarity0_r = interface4_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank4_ev_polarity0_we <= 1'd0;
    csrbank4_ev_polarity0_re <= 1'd0;
    if ((csrbank4_sel & (interface4_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank4_ev_polarity0_re <= interface4_bank_bus_we;
        csrbank4_ev_polarity0_we <= csrbank4_re;
    end
end
assign csrbank4_ev_status_r = interface4_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank4_ev_status_re <= 1'd0;
    csrbank4_ev_status_we <= 1'd0;
    if ((csrbank4_sel & (interface4_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank4_ev_status_re <= interface4_bank_bus_we;
        csrbank4_ev_status_we <= csrbank4_re;
    end
end
assign csrbank4_ev_pending_r = interface4_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank4_ev_pending_we <= 1'd0;
    csrbank4_ev_pending_re <= 1'd0;
    if ((csrbank4_sel & (interface4_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank4_ev_pending_re <= interface4_bank_bus_we;
        csrbank4_ev_pending_we <= csrbank4_re;
    end
end
assign csrbank4_ev_enable0_r = interface4_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank4_ev_enable0_we <= 1'd0;
    csrbank4_ev_enable0_re <= 1'd0;
    if ((csrbank4_sel & (interface4_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank4_ev_enable0_re <= interface4_bank_bus_we;
        csrbank4_ev_enable0_we <= csrbank4_re;
    end
end
always @(*) begin
    irqarray1_trigger <= 16'd0;
    if (irqarray1_soft_re) begin
        irqarray1_trigger <= irqarray1_soft_storage[15:0];
    end
end
assign csrbank4_ev_soft0_w = irqarray1_soft_storage[15:0];
assign irqarray1_use_edge = irqarray1_edge_triggered_storage[15:0];
assign csrbank4_ev_edge_triggered0_w = irqarray1_edge_triggered_storage[15:0];
assign irqarray1_rising = irqarray1_polarity_storage[15:0];
assign csrbank4_ev_polarity0_w = irqarray1_polarity_storage[15:0];
always @(*) begin
    irqarray1_status_status <= 16'd0;
    irqarray1_status_status[0] <= irqarray1_usbc_dupe0;
    irqarray1_status_status[1] <= irqarray1_nc_b1s10;
    irqarray1_status_status[2] <= irqarray1_nc_b1s20;
    irqarray1_status_status[3] <= irqarray1_nc_b1s30;
    irqarray1_status_status[4] <= irqarray1_nc_b1s40;
    irqarray1_status_status[5] <= irqarray1_nc_b1s50;
    irqarray1_status_status[6] <= irqarray1_nc_b1s60;
    irqarray1_status_status[7] <= irqarray1_nc_b1s70;
    irqarray1_status_status[8] <= irqarray1_nc_b1s80;
    irqarray1_status_status[9] <= irqarray1_nc_b1s90;
    irqarray1_status_status[10] <= irqarray1_nc_b1s100;
    irqarray1_status_status[11] <= irqarray1_nc_b1s110;
    irqarray1_status_status[12] <= irqarray1_nc_b1s120;
    irqarray1_status_status[13] <= irqarray1_nc_b1s130;
    irqarray1_status_status[14] <= irqarray1_nc_b1s140;
    irqarray1_status_status[15] <= irqarray1_nc_b1s150;
end
assign csrbank4_ev_status_w = irqarray1_status_status[15:0];
assign irqarray1_status_we = csrbank4_ev_status_we;
always @(*) begin
    irqarray1_pending_status <= 16'd0;
    irqarray1_pending_status[0] <= irqarray1_usbc_dupe1;
    irqarray1_pending_status[1] <= irqarray1_nc_b1s11;
    irqarray1_pending_status[2] <= irqarray1_nc_b1s21;
    irqarray1_pending_status[3] <= irqarray1_nc_b1s31;
    irqarray1_pending_status[4] <= irqarray1_nc_b1s41;
    irqarray1_pending_status[5] <= irqarray1_nc_b1s51;
    irqarray1_pending_status[6] <= irqarray1_nc_b1s61;
    irqarray1_pending_status[7] <= irqarray1_nc_b1s71;
    irqarray1_pending_status[8] <= irqarray1_nc_b1s81;
    irqarray1_pending_status[9] <= irqarray1_nc_b1s91;
    irqarray1_pending_status[10] <= irqarray1_nc_b1s101;
    irqarray1_pending_status[11] <= irqarray1_nc_b1s111;
    irqarray1_pending_status[12] <= irqarray1_nc_b1s121;
    irqarray1_pending_status[13] <= irqarray1_nc_b1s131;
    irqarray1_pending_status[14] <= irqarray1_nc_b1s141;
    irqarray1_pending_status[15] <= irqarray1_nc_b1s151;
end
assign csrbank4_ev_pending_w = irqarray1_pending_status[15:0];
assign irqarray1_pending_we = csrbank4_ev_pending_we;
assign irqarray1_usbc_dupe2 = irqarray1_enable_storage[0];
assign irqarray1_nc_b1s12 = irqarray1_enable_storage[1];
assign irqarray1_nc_b1s22 = irqarray1_enable_storage[2];
assign irqarray1_nc_b1s32 = irqarray1_enable_storage[3];
assign irqarray1_nc_b1s42 = irqarray1_enable_storage[4];
assign irqarray1_nc_b1s52 = irqarray1_enable_storage[5];
assign irqarray1_nc_b1s62 = irqarray1_enable_storage[6];
assign irqarray1_nc_b1s72 = irqarray1_enable_storage[7];
assign irqarray1_nc_b1s82 = irqarray1_enable_storage[8];
assign irqarray1_nc_b1s92 = irqarray1_enable_storage[9];
assign irqarray1_nc_b1s102 = irqarray1_enable_storage[10];
assign irqarray1_nc_b1s112 = irqarray1_enable_storage[11];
assign irqarray1_nc_b1s122 = irqarray1_enable_storage[12];
assign irqarray1_nc_b1s132 = irqarray1_enable_storage[13];
assign irqarray1_nc_b1s142 = irqarray1_enable_storage[14];
assign irqarray1_nc_b1s152 = irqarray1_enable_storage[15];
assign csrbank4_ev_enable0_w = irqarray1_enable_storage[15:0];
assign csrbank5_sel = (interface5_bank_bus_adr[15:10] == 3'd6);
assign csrbank5_re = interface5_bank_bus_re;
assign csrbank5_ev_soft0_r = interface5_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank5_ev_soft0_re <= 1'd0;
    csrbank5_ev_soft0_we <= 1'd0;
    if ((csrbank5_sel & (interface5_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank5_ev_soft0_re <= interface5_bank_bus_we;
        csrbank5_ev_soft0_we <= csrbank5_re;
    end
end
assign csrbank5_ev_edge_triggered0_r = interface5_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank5_ev_edge_triggered0_we <= 1'd0;
    csrbank5_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank5_sel & (interface5_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank5_ev_edge_triggered0_re <= interface5_bank_bus_we;
        csrbank5_ev_edge_triggered0_we <= csrbank5_re;
    end
end
assign csrbank5_ev_polarity0_r = interface5_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank5_ev_polarity0_we <= 1'd0;
    csrbank5_ev_polarity0_re <= 1'd0;
    if ((csrbank5_sel & (interface5_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank5_ev_polarity0_re <= interface5_bank_bus_we;
        csrbank5_ev_polarity0_we <= csrbank5_re;
    end
end
assign csrbank5_ev_status_r = interface5_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank5_ev_status_re <= 1'd0;
    csrbank5_ev_status_we <= 1'd0;
    if ((csrbank5_sel & (interface5_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank5_ev_status_re <= interface5_bank_bus_we;
        csrbank5_ev_status_we <= csrbank5_re;
    end
end
assign csrbank5_ev_pending_r = interface5_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank5_ev_pending_we <= 1'd0;
    csrbank5_ev_pending_re <= 1'd0;
    if ((csrbank5_sel & (interface5_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank5_ev_pending_re <= interface5_bank_bus_we;
        csrbank5_ev_pending_we <= csrbank5_re;
    end
end
assign csrbank5_ev_enable0_r = interface5_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank5_ev_enable0_we <= 1'd0;
    csrbank5_ev_enable0_re <= 1'd0;
    if ((csrbank5_sel & (interface5_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank5_ev_enable0_re <= interface5_bank_bus_we;
        csrbank5_ev_enable0_we <= csrbank5_re;
    end
end
always @(*) begin
    irqarray10_trigger <= 16'd0;
    if (irqarray10_soft_re) begin
        irqarray10_trigger <= irqarray10_soft_storage[15:0];
    end
end
assign csrbank5_ev_soft0_w = irqarray10_soft_storage[15:0];
assign irqarray10_use_edge = irqarray10_edge_triggered_storage[15:0];
assign csrbank5_ev_edge_triggered0_w = irqarray10_edge_triggered_storage[15:0];
assign irqarray10_rising = irqarray10_polarity_storage[15:0];
assign csrbank5_ev_polarity0_w = irqarray10_polarity_storage[15:0];
always @(*) begin
    irqarray10_status_status <= 16'd0;
    irqarray10_status_status[0] <= irqarray10_ioxirq0;
    irqarray10_status_status[1] <= irqarray10_usbc0;
    irqarray10_status_status[2] <= irqarray10_sddcirq0;
    irqarray10_status_status[3] <= irqarray10_pioirq00;
    irqarray10_status_status[4] <= irqarray10_pioirq10;
    irqarray10_status_status[5] <= irqarray10_pioirq20;
    irqarray10_status_status[6] <= irqarray10_pioirq30;
    irqarray10_status_status[7] <= irqarray10_nc_b10s70;
    irqarray10_status_status[8] <= irqarray10_nc_b10s80;
    irqarray10_status_status[9] <= irqarray10_nc_b10s90;
    irqarray10_status_status[10] <= irqarray10_nc_b10s100;
    irqarray10_status_status[11] <= irqarray10_nc_b10s110;
    irqarray10_status_status[12] <= irqarray10_nc_b10s120;
    irqarray10_status_status[13] <= irqarray10_nc_b10s130;
    irqarray10_status_status[14] <= irqarray10_nc_b10s140;
    irqarray10_status_status[15] <= irqarray10_nc_b10s150;
end
assign csrbank5_ev_status_w = irqarray10_status_status[15:0];
assign irqarray10_status_we = csrbank5_ev_status_we;
always @(*) begin
    irqarray10_pending_status <= 16'd0;
    irqarray10_pending_status[0] <= irqarray10_ioxirq1;
    irqarray10_pending_status[1] <= irqarray10_usbc1;
    irqarray10_pending_status[2] <= irqarray10_sddcirq1;
    irqarray10_pending_status[3] <= irqarray10_pioirq01;
    irqarray10_pending_status[4] <= irqarray10_pioirq11;
    irqarray10_pending_status[5] <= irqarray10_pioirq21;
    irqarray10_pending_status[6] <= irqarray10_pioirq31;
    irqarray10_pending_status[7] <= irqarray10_nc_b10s71;
    irqarray10_pending_status[8] <= irqarray10_nc_b10s81;
    irqarray10_pending_status[9] <= irqarray10_nc_b10s91;
    irqarray10_pending_status[10] <= irqarray10_nc_b10s101;
    irqarray10_pending_status[11] <= irqarray10_nc_b10s111;
    irqarray10_pending_status[12] <= irqarray10_nc_b10s121;
    irqarray10_pending_status[13] <= irqarray10_nc_b10s131;
    irqarray10_pending_status[14] <= irqarray10_nc_b10s141;
    irqarray10_pending_status[15] <= irqarray10_nc_b10s151;
end
assign csrbank5_ev_pending_w = irqarray10_pending_status[15:0];
assign irqarray10_pending_we = csrbank5_ev_pending_we;
assign irqarray10_ioxirq2 = irqarray10_enable_storage[0];
assign irqarray10_usbc2 = irqarray10_enable_storage[1];
assign irqarray10_sddcirq2 = irqarray10_enable_storage[2];
assign irqarray10_pioirq02 = irqarray10_enable_storage[3];
assign irqarray10_pioirq12 = irqarray10_enable_storage[4];
assign irqarray10_pioirq22 = irqarray10_enable_storage[5];
assign irqarray10_pioirq32 = irqarray10_enable_storage[6];
assign irqarray10_nc_b10s72 = irqarray10_enable_storage[7];
assign irqarray10_nc_b10s82 = irqarray10_enable_storage[8];
assign irqarray10_nc_b10s92 = irqarray10_enable_storage[9];
assign irqarray10_nc_b10s102 = irqarray10_enable_storage[10];
assign irqarray10_nc_b10s112 = irqarray10_enable_storage[11];
assign irqarray10_nc_b10s122 = irqarray10_enable_storage[12];
assign irqarray10_nc_b10s132 = irqarray10_enable_storage[13];
assign irqarray10_nc_b10s142 = irqarray10_enable_storage[14];
assign irqarray10_nc_b10s152 = irqarray10_enable_storage[15];
assign csrbank5_ev_enable0_w = irqarray10_enable_storage[15:0];
assign csrbank6_sel = (interface6_bank_bus_adr[15:10] == 3'd7);
assign csrbank6_re = interface6_bank_bus_re;
assign csrbank6_ev_soft0_r = interface6_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank6_ev_soft0_re <= 1'd0;
    csrbank6_ev_soft0_we <= 1'd0;
    if ((csrbank6_sel & (interface6_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank6_ev_soft0_re <= interface6_bank_bus_we;
        csrbank6_ev_soft0_we <= csrbank6_re;
    end
end
assign csrbank6_ev_edge_triggered0_r = interface6_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank6_ev_edge_triggered0_we <= 1'd0;
    csrbank6_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank6_sel & (interface6_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank6_ev_edge_triggered0_re <= interface6_bank_bus_we;
        csrbank6_ev_edge_triggered0_we <= csrbank6_re;
    end
end
assign csrbank6_ev_polarity0_r = interface6_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank6_ev_polarity0_we <= 1'd0;
    csrbank6_ev_polarity0_re <= 1'd0;
    if ((csrbank6_sel & (interface6_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank6_ev_polarity0_re <= interface6_bank_bus_we;
        csrbank6_ev_polarity0_we <= csrbank6_re;
    end
end
assign csrbank6_ev_status_r = interface6_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank6_ev_status_re <= 1'd0;
    csrbank6_ev_status_we <= 1'd0;
    if ((csrbank6_sel & (interface6_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank6_ev_status_re <= interface6_bank_bus_we;
        csrbank6_ev_status_we <= csrbank6_re;
    end
end
assign csrbank6_ev_pending_r = interface6_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank6_ev_pending_we <= 1'd0;
    csrbank6_ev_pending_re <= 1'd0;
    if ((csrbank6_sel & (interface6_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank6_ev_pending_re <= interface6_bank_bus_we;
        csrbank6_ev_pending_we <= csrbank6_re;
    end
end
assign csrbank6_ev_enable0_r = interface6_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank6_ev_enable0_we <= 1'd0;
    csrbank6_ev_enable0_re <= 1'd0;
    if ((csrbank6_sel & (interface6_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank6_ev_enable0_re <= interface6_bank_bus_we;
        csrbank6_ev_enable0_we <= csrbank6_re;
    end
end
always @(*) begin
    irqarray11_trigger <= 16'd0;
    if (irqarray11_soft_re) begin
        irqarray11_trigger <= irqarray11_soft_storage[15:0];
    end
end
assign csrbank6_ev_soft0_w = irqarray11_soft_storage[15:0];
assign irqarray11_use_edge = irqarray11_edge_triggered_storage[15:0];
assign csrbank6_ev_edge_triggered0_w = irqarray11_edge_triggered_storage[15:0];
assign irqarray11_rising = irqarray11_polarity_storage[15:0];
assign csrbank6_ev_polarity0_w = irqarray11_polarity_storage[15:0];
always @(*) begin
    irqarray11_status_status <= 16'd0;
    irqarray11_status_status[0] <= irqarray11_i2s_rx_dupe0;
    irqarray11_status_status[1] <= irqarray11_i2s_tx_dupe0;
    irqarray11_status_status[2] <= irqarray11_nc_b11s20;
    irqarray11_status_status[3] <= irqarray11_nc_b11s30;
    irqarray11_status_status[4] <= irqarray11_nc_b11s40;
    irqarray11_status_status[5] <= irqarray11_nc_b11s50;
    irqarray11_status_status[6] <= irqarray11_nc_b11s60;
    irqarray11_status_status[7] <= irqarray11_nc_b11s70;
    irqarray11_status_status[8] <= irqarray11_nc_b11s80;
    irqarray11_status_status[9] <= irqarray11_nc_b11s90;
    irqarray11_status_status[10] <= irqarray11_nc_b11s100;
    irqarray11_status_status[11] <= irqarray11_nc_b11s110;
    irqarray11_status_status[12] <= irqarray11_nc_b11s120;
    irqarray11_status_status[13] <= irqarray11_nc_b11s130;
    irqarray11_status_status[14] <= irqarray11_nc_b11s140;
    irqarray11_status_status[15] <= irqarray11_nc_b11s150;
end
assign csrbank6_ev_status_w = irqarray11_status_status[15:0];
assign irqarray11_status_we = csrbank6_ev_status_we;
always @(*) begin
    irqarray11_pending_status <= 16'd0;
    irqarray11_pending_status[0] <= irqarray11_i2s_rx_dupe1;
    irqarray11_pending_status[1] <= irqarray11_i2s_tx_dupe1;
    irqarray11_pending_status[2] <= irqarray11_nc_b11s21;
    irqarray11_pending_status[3] <= irqarray11_nc_b11s31;
    irqarray11_pending_status[4] <= irqarray11_nc_b11s41;
    irqarray11_pending_status[5] <= irqarray11_nc_b11s51;
    irqarray11_pending_status[6] <= irqarray11_nc_b11s61;
    irqarray11_pending_status[7] <= irqarray11_nc_b11s71;
    irqarray11_pending_status[8] <= irqarray11_nc_b11s81;
    irqarray11_pending_status[9] <= irqarray11_nc_b11s91;
    irqarray11_pending_status[10] <= irqarray11_nc_b11s101;
    irqarray11_pending_status[11] <= irqarray11_nc_b11s111;
    irqarray11_pending_status[12] <= irqarray11_nc_b11s121;
    irqarray11_pending_status[13] <= irqarray11_nc_b11s131;
    irqarray11_pending_status[14] <= irqarray11_nc_b11s141;
    irqarray11_pending_status[15] <= irqarray11_nc_b11s151;
end
assign csrbank6_ev_pending_w = irqarray11_pending_status[15:0];
assign irqarray11_pending_we = csrbank6_ev_pending_we;
assign irqarray11_i2s_rx_dupe2 = irqarray11_enable_storage[0];
assign irqarray11_i2s_tx_dupe2 = irqarray11_enable_storage[1];
assign irqarray11_nc_b11s22 = irqarray11_enable_storage[2];
assign irqarray11_nc_b11s32 = irqarray11_enable_storage[3];
assign irqarray11_nc_b11s42 = irqarray11_enable_storage[4];
assign irqarray11_nc_b11s52 = irqarray11_enable_storage[5];
assign irqarray11_nc_b11s62 = irqarray11_enable_storage[6];
assign irqarray11_nc_b11s72 = irqarray11_enable_storage[7];
assign irqarray11_nc_b11s82 = irqarray11_enable_storage[8];
assign irqarray11_nc_b11s92 = irqarray11_enable_storage[9];
assign irqarray11_nc_b11s102 = irqarray11_enable_storage[10];
assign irqarray11_nc_b11s112 = irqarray11_enable_storage[11];
assign irqarray11_nc_b11s122 = irqarray11_enable_storage[12];
assign irqarray11_nc_b11s132 = irqarray11_enable_storage[13];
assign irqarray11_nc_b11s142 = irqarray11_enable_storage[14];
assign irqarray11_nc_b11s152 = irqarray11_enable_storage[15];
assign csrbank6_ev_enable0_w = irqarray11_enable_storage[15:0];
assign csrbank7_sel = (interface7_bank_bus_adr[15:10] == 4'd8);
assign csrbank7_re = interface7_bank_bus_re;
assign csrbank7_ev_soft0_r = interface7_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank7_ev_soft0_re <= 1'd0;
    csrbank7_ev_soft0_we <= 1'd0;
    if ((csrbank7_sel & (interface7_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank7_ev_soft0_re <= interface7_bank_bus_we;
        csrbank7_ev_soft0_we <= csrbank7_re;
    end
end
assign csrbank7_ev_edge_triggered0_r = interface7_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank7_ev_edge_triggered0_we <= 1'd0;
    csrbank7_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank7_sel & (interface7_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank7_ev_edge_triggered0_re <= interface7_bank_bus_we;
        csrbank7_ev_edge_triggered0_we <= csrbank7_re;
    end
end
assign csrbank7_ev_polarity0_r = interface7_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank7_ev_polarity0_we <= 1'd0;
    csrbank7_ev_polarity0_re <= 1'd0;
    if ((csrbank7_sel & (interface7_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank7_ev_polarity0_re <= interface7_bank_bus_we;
        csrbank7_ev_polarity0_we <= csrbank7_re;
    end
end
assign csrbank7_ev_status_r = interface7_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank7_ev_status_re <= 1'd0;
    csrbank7_ev_status_we <= 1'd0;
    if ((csrbank7_sel & (interface7_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank7_ev_status_re <= interface7_bank_bus_we;
        csrbank7_ev_status_we <= csrbank7_re;
    end
end
assign csrbank7_ev_pending_r = interface7_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank7_ev_pending_we <= 1'd0;
    csrbank7_ev_pending_re <= 1'd0;
    if ((csrbank7_sel & (interface7_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank7_ev_pending_re <= interface7_bank_bus_we;
        csrbank7_ev_pending_we <= csrbank7_re;
    end
end
assign csrbank7_ev_enable0_r = interface7_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank7_ev_enable0_we <= 1'd0;
    csrbank7_ev_enable0_re <= 1'd0;
    if ((csrbank7_sel & (interface7_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank7_ev_enable0_re <= interface7_bank_bus_we;
        csrbank7_ev_enable0_we <= csrbank7_re;
    end
end
always @(*) begin
    irqarray12_trigger <= 16'd0;
    if (irqarray12_soft_re) begin
        irqarray12_trigger <= irqarray12_soft_storage[15:0];
    end
end
assign csrbank7_ev_soft0_w = irqarray12_soft_storage[15:0];
assign irqarray12_use_edge = irqarray12_edge_triggered_storage[15:0];
assign csrbank7_ev_edge_triggered0_w = irqarray12_edge_triggered_storage[15:0];
assign irqarray12_rising = irqarray12_polarity_storage[15:0];
assign csrbank7_ev_polarity0_w = irqarray12_polarity_storage[15:0];
always @(*) begin
    irqarray12_status_status <= 16'd0;
    irqarray12_status_status[0] <= irqarray12_nc_b12s00;
    irqarray12_status_status[1] <= irqarray12_nc_b12s10;
    irqarray12_status_status[2] <= irqarray12_nc_b12s20;
    irqarray12_status_status[3] <= irqarray12_nc_b12s30;
    irqarray12_status_status[4] <= irqarray12_nc_b12s40;
    irqarray12_status_status[5] <= irqarray12_nc_b12s50;
    irqarray12_status_status[6] <= irqarray12_nc_b12s60;
    irqarray12_status_status[7] <= irqarray12_nc_b12s70;
    irqarray12_status_status[8] <= irqarray12_i2c0_nack0;
    irqarray12_status_status[9] <= irqarray12_i2c1_nack0;
    irqarray12_status_status[10] <= irqarray12_i2c2_nack0;
    irqarray12_status_status[11] <= irqarray12_i2c3_nack0;
    irqarray12_status_status[12] <= irqarray12_i2c0_err0;
    irqarray12_status_status[13] <= irqarray12_i2c1_err0;
    irqarray12_status_status[14] <= irqarray12_i2c2_err0;
    irqarray12_status_status[15] <= irqarray12_i2c3_err0;
end
assign csrbank7_ev_status_w = irqarray12_status_status[15:0];
assign irqarray12_status_we = csrbank7_ev_status_we;
always @(*) begin
    irqarray12_pending_status <= 16'd0;
    irqarray12_pending_status[0] <= irqarray12_nc_b12s01;
    irqarray12_pending_status[1] <= irqarray12_nc_b12s11;
    irqarray12_pending_status[2] <= irqarray12_nc_b12s21;
    irqarray12_pending_status[3] <= irqarray12_nc_b12s31;
    irqarray12_pending_status[4] <= irqarray12_nc_b12s41;
    irqarray12_pending_status[5] <= irqarray12_nc_b12s51;
    irqarray12_pending_status[6] <= irqarray12_nc_b12s61;
    irqarray12_pending_status[7] <= irqarray12_nc_b12s71;
    irqarray12_pending_status[8] <= irqarray12_i2c0_nack1;
    irqarray12_pending_status[9] <= irqarray12_i2c1_nack1;
    irqarray12_pending_status[10] <= irqarray12_i2c2_nack1;
    irqarray12_pending_status[11] <= irqarray12_i2c3_nack1;
    irqarray12_pending_status[12] <= irqarray12_i2c0_err1;
    irqarray12_pending_status[13] <= irqarray12_i2c1_err1;
    irqarray12_pending_status[14] <= irqarray12_i2c2_err1;
    irqarray12_pending_status[15] <= irqarray12_i2c3_err1;
end
assign csrbank7_ev_pending_w = irqarray12_pending_status[15:0];
assign irqarray12_pending_we = csrbank7_ev_pending_we;
assign irqarray12_nc_b12s02 = irqarray12_enable_storage[0];
assign irqarray12_nc_b12s12 = irqarray12_enable_storage[1];
assign irqarray12_nc_b12s22 = irqarray12_enable_storage[2];
assign irqarray12_nc_b12s32 = irqarray12_enable_storage[3];
assign irqarray12_nc_b12s42 = irqarray12_enable_storage[4];
assign irqarray12_nc_b12s52 = irqarray12_enable_storage[5];
assign irqarray12_nc_b12s62 = irqarray12_enable_storage[6];
assign irqarray12_nc_b12s72 = irqarray12_enable_storage[7];
assign irqarray12_i2c0_nack2 = irqarray12_enable_storage[8];
assign irqarray12_i2c1_nack2 = irqarray12_enable_storage[9];
assign irqarray12_i2c2_nack2 = irqarray12_enable_storage[10];
assign irqarray12_i2c3_nack2 = irqarray12_enable_storage[11];
assign irqarray12_i2c0_err2 = irqarray12_enable_storage[12];
assign irqarray12_i2c1_err2 = irqarray12_enable_storage[13];
assign irqarray12_i2c2_err2 = irqarray12_enable_storage[14];
assign irqarray12_i2c3_err2 = irqarray12_enable_storage[15];
assign csrbank7_ev_enable0_w = irqarray12_enable_storage[15:0];
assign csrbank8_sel = (interface8_bank_bus_adr[15:10] == 4'd9);
assign csrbank8_re = interface8_bank_bus_re;
assign csrbank8_ev_soft0_r = interface8_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank8_ev_soft0_re <= 1'd0;
    csrbank8_ev_soft0_we <= 1'd0;
    if ((csrbank8_sel & (interface8_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank8_ev_soft0_re <= interface8_bank_bus_we;
        csrbank8_ev_soft0_we <= csrbank8_re;
    end
end
assign csrbank8_ev_edge_triggered0_r = interface8_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank8_ev_edge_triggered0_we <= 1'd0;
    csrbank8_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank8_sel & (interface8_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank8_ev_edge_triggered0_re <= interface8_bank_bus_we;
        csrbank8_ev_edge_triggered0_we <= csrbank8_re;
    end
end
assign csrbank8_ev_polarity0_r = interface8_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank8_ev_polarity0_we <= 1'd0;
    csrbank8_ev_polarity0_re <= 1'd0;
    if ((csrbank8_sel & (interface8_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank8_ev_polarity0_re <= interface8_bank_bus_we;
        csrbank8_ev_polarity0_we <= csrbank8_re;
    end
end
assign csrbank8_ev_status_r = interface8_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank8_ev_status_re <= 1'd0;
    csrbank8_ev_status_we <= 1'd0;
    if ((csrbank8_sel & (interface8_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank8_ev_status_re <= interface8_bank_bus_we;
        csrbank8_ev_status_we <= csrbank8_re;
    end
end
assign csrbank8_ev_pending_r = interface8_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank8_ev_pending_we <= 1'd0;
    csrbank8_ev_pending_re <= 1'd0;
    if ((csrbank8_sel & (interface8_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank8_ev_pending_re <= interface8_bank_bus_we;
        csrbank8_ev_pending_we <= csrbank8_re;
    end
end
assign csrbank8_ev_enable0_r = interface8_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank8_ev_enable0_we <= 1'd0;
    csrbank8_ev_enable0_re <= 1'd0;
    if ((csrbank8_sel & (interface8_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank8_ev_enable0_re <= interface8_bank_bus_we;
        csrbank8_ev_enable0_we <= csrbank8_re;
    end
end
always @(*) begin
    irqarray13_trigger <= 16'd0;
    if (irqarray13_soft_re) begin
        irqarray13_trigger <= irqarray13_soft_storage[15:0];
    end
end
assign csrbank8_ev_soft0_w = irqarray13_soft_storage[15:0];
assign irqarray13_use_edge = irqarray13_edge_triggered_storage[15:0];
assign csrbank8_ev_edge_triggered0_w = irqarray13_edge_triggered_storage[15:0];
assign irqarray13_rising = irqarray13_polarity_storage[15:0];
assign csrbank8_ev_polarity0_w = irqarray13_polarity_storage[15:0];
always @(*) begin
    irqarray13_status_status <= 16'd0;
    irqarray13_status_status[0] <= irqarray13_coresuberr0;
    irqarray13_status_status[1] <= irqarray13_sceerr0;
    irqarray13_status_status[2] <= irqarray13_ifsuberr0;
    irqarray13_status_status[3] <= irqarray13_secirq0;
    irqarray13_status_status[4] <= irqarray13_nc_b13s40;
    irqarray13_status_status[5] <= irqarray13_nc_b13s50;
    irqarray13_status_status[6] <= irqarray13_nc_b13s60;
    irqarray13_status_status[7] <= irqarray13_nc_b13s70;
    irqarray13_status_status[8] <= irqarray13_nc_b13s80;
    irqarray13_status_status[9] <= irqarray13_nc_b13s90;
    irqarray13_status_status[10] <= irqarray13_nc_b13s100;
    irqarray13_status_status[11] <= irqarray13_nc_b13s110;
    irqarray13_status_status[12] <= irqarray13_nc_b13s120;
    irqarray13_status_status[13] <= irqarray13_nc_b13s130;
    irqarray13_status_status[14] <= irqarray13_nc_b13s140;
    irqarray13_status_status[15] <= irqarray13_nc_b13s150;
end
assign csrbank8_ev_status_w = irqarray13_status_status[15:0];
assign irqarray13_status_we = csrbank8_ev_status_we;
always @(*) begin
    irqarray13_pending_status <= 16'd0;
    irqarray13_pending_status[0] <= irqarray13_coresuberr1;
    irqarray13_pending_status[1] <= irqarray13_sceerr1;
    irqarray13_pending_status[2] <= irqarray13_ifsuberr1;
    irqarray13_pending_status[3] <= irqarray13_secirq1;
    irqarray13_pending_status[4] <= irqarray13_nc_b13s41;
    irqarray13_pending_status[5] <= irqarray13_nc_b13s51;
    irqarray13_pending_status[6] <= irqarray13_nc_b13s61;
    irqarray13_pending_status[7] <= irqarray13_nc_b13s71;
    irqarray13_pending_status[8] <= irqarray13_nc_b13s81;
    irqarray13_pending_status[9] <= irqarray13_nc_b13s91;
    irqarray13_pending_status[10] <= irqarray13_nc_b13s101;
    irqarray13_pending_status[11] <= irqarray13_nc_b13s111;
    irqarray13_pending_status[12] <= irqarray13_nc_b13s121;
    irqarray13_pending_status[13] <= irqarray13_nc_b13s131;
    irqarray13_pending_status[14] <= irqarray13_nc_b13s141;
    irqarray13_pending_status[15] <= irqarray13_nc_b13s151;
end
assign csrbank8_ev_pending_w = irqarray13_pending_status[15:0];
assign irqarray13_pending_we = csrbank8_ev_pending_we;
assign irqarray13_coresuberr2 = irqarray13_enable_storage[0];
assign irqarray13_sceerr2 = irqarray13_enable_storage[1];
assign irqarray13_ifsuberr2 = irqarray13_enable_storage[2];
assign irqarray13_secirq2 = irqarray13_enable_storage[3];
assign irqarray13_nc_b13s42 = irqarray13_enable_storage[4];
assign irqarray13_nc_b13s52 = irqarray13_enable_storage[5];
assign irqarray13_nc_b13s62 = irqarray13_enable_storage[6];
assign irqarray13_nc_b13s72 = irqarray13_enable_storage[7];
assign irqarray13_nc_b13s82 = irqarray13_enable_storage[8];
assign irqarray13_nc_b13s92 = irqarray13_enable_storage[9];
assign irqarray13_nc_b13s102 = irqarray13_enable_storage[10];
assign irqarray13_nc_b13s112 = irqarray13_enable_storage[11];
assign irqarray13_nc_b13s122 = irqarray13_enable_storage[12];
assign irqarray13_nc_b13s132 = irqarray13_enable_storage[13];
assign irqarray13_nc_b13s142 = irqarray13_enable_storage[14];
assign irqarray13_nc_b13s152 = irqarray13_enable_storage[15];
assign csrbank8_ev_enable0_w = irqarray13_enable_storage[15:0];
assign csrbank9_sel = (interface9_bank_bus_adr[15:10] == 4'd10);
assign csrbank9_re = interface9_bank_bus_re;
assign csrbank9_ev_soft0_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank9_ev_soft0_re <= 1'd0;
    csrbank9_ev_soft0_we <= 1'd0;
    if ((csrbank9_sel & (interface9_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank9_ev_soft0_re <= interface9_bank_bus_we;
        csrbank9_ev_soft0_we <= csrbank9_re;
    end
end
assign csrbank9_ev_edge_triggered0_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank9_ev_edge_triggered0_we <= 1'd0;
    csrbank9_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank9_sel & (interface9_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank9_ev_edge_triggered0_re <= interface9_bank_bus_we;
        csrbank9_ev_edge_triggered0_we <= csrbank9_re;
    end
end
assign csrbank9_ev_polarity0_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank9_ev_polarity0_we <= 1'd0;
    csrbank9_ev_polarity0_re <= 1'd0;
    if ((csrbank9_sel & (interface9_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank9_ev_polarity0_re <= interface9_bank_bus_we;
        csrbank9_ev_polarity0_we <= csrbank9_re;
    end
end
assign csrbank9_ev_status_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank9_ev_status_re <= 1'd0;
    csrbank9_ev_status_we <= 1'd0;
    if ((csrbank9_sel & (interface9_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank9_ev_status_re <= interface9_bank_bus_we;
        csrbank9_ev_status_we <= csrbank9_re;
    end
end
assign csrbank9_ev_pending_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank9_ev_pending_we <= 1'd0;
    csrbank9_ev_pending_re <= 1'd0;
    if ((csrbank9_sel & (interface9_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank9_ev_pending_re <= interface9_bank_bus_we;
        csrbank9_ev_pending_we <= csrbank9_re;
    end
end
assign csrbank9_ev_enable0_r = interface9_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank9_ev_enable0_we <= 1'd0;
    csrbank9_ev_enable0_re <= 1'd0;
    if ((csrbank9_sel & (interface9_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank9_ev_enable0_re <= interface9_bank_bus_we;
        csrbank9_ev_enable0_we <= csrbank9_re;
    end
end
always @(*) begin
    irqarray14_trigger <= 16'd0;
    if (irqarray14_soft_re) begin
        irqarray14_trigger <= irqarray14_soft_storage[15:0];
    end
end
assign csrbank9_ev_soft0_w = irqarray14_soft_storage[15:0];
assign irqarray14_use_edge = irqarray14_edge_triggered_storage[15:0];
assign csrbank9_ev_edge_triggered0_w = irqarray14_edge_triggered_storage[15:0];
assign irqarray14_rising = irqarray14_polarity_storage[15:0];
assign csrbank9_ev_polarity0_w = irqarray14_polarity_storage[15:0];
always @(*) begin
    irqarray14_status_status <= 16'd0;
    irqarray14_status_status[0] <= irqarray14_uart2_rx_dupe0;
    irqarray14_status_status[1] <= irqarray14_uart2_tx_dupe0;
    irqarray14_status_status[2] <= irqarray14_uart2_rx_char_dupe0;
    irqarray14_status_status[3] <= irqarray14_uart2_err_dupe0;
    irqarray14_status_status[4] <= irqarray14_uart3_rx_dupe0;
    irqarray14_status_status[5] <= irqarray14_uart3_tx_dupe0;
    irqarray14_status_status[6] <= irqarray14_uart3_rx_char_dupe0;
    irqarray14_status_status[7] <= irqarray14_uart3_err_dupe0;
    irqarray14_status_status[8] <= irqarray14_trng_done_dupe0;
    irqarray14_status_status[9] <= irqarray14_nc_b14s90;
    irqarray14_status_status[10] <= irqarray14_nc_b14s100;
    irqarray14_status_status[11] <= irqarray14_nc_b14s110;
    irqarray14_status_status[12] <= irqarray14_nc_b14s120;
    irqarray14_status_status[13] <= irqarray14_nc_b14s130;
    irqarray14_status_status[14] <= irqarray14_nc_b14s140;
    irqarray14_status_status[15] <= irqarray14_nc_b14s150;
end
assign csrbank9_ev_status_w = irqarray14_status_status[15:0];
assign irqarray14_status_we = csrbank9_ev_status_we;
always @(*) begin
    irqarray14_pending_status <= 16'd0;
    irqarray14_pending_status[0] <= irqarray14_uart2_rx_dupe1;
    irqarray14_pending_status[1] <= irqarray14_uart2_tx_dupe1;
    irqarray14_pending_status[2] <= irqarray14_uart2_rx_char_dupe1;
    irqarray14_pending_status[3] <= irqarray14_uart2_err_dupe1;
    irqarray14_pending_status[4] <= irqarray14_uart3_rx_dupe1;
    irqarray14_pending_status[5] <= irqarray14_uart3_tx_dupe1;
    irqarray14_pending_status[6] <= irqarray14_uart3_rx_char_dupe1;
    irqarray14_pending_status[7] <= irqarray14_uart3_err_dupe1;
    irqarray14_pending_status[8] <= irqarray14_trng_done_dupe1;
    irqarray14_pending_status[9] <= irqarray14_nc_b14s91;
    irqarray14_pending_status[10] <= irqarray14_nc_b14s101;
    irqarray14_pending_status[11] <= irqarray14_nc_b14s111;
    irqarray14_pending_status[12] <= irqarray14_nc_b14s121;
    irqarray14_pending_status[13] <= irqarray14_nc_b14s131;
    irqarray14_pending_status[14] <= irqarray14_nc_b14s141;
    irqarray14_pending_status[15] <= irqarray14_nc_b14s151;
end
assign csrbank9_ev_pending_w = irqarray14_pending_status[15:0];
assign irqarray14_pending_we = csrbank9_ev_pending_we;
assign irqarray14_uart2_rx_dupe2 = irqarray14_enable_storage[0];
assign irqarray14_uart2_tx_dupe2 = irqarray14_enable_storage[1];
assign irqarray14_uart2_rx_char_dupe2 = irqarray14_enable_storage[2];
assign irqarray14_uart2_err_dupe2 = irqarray14_enable_storage[3];
assign irqarray14_uart3_rx_dupe2 = irqarray14_enable_storage[4];
assign irqarray14_uart3_tx_dupe2 = irqarray14_enable_storage[5];
assign irqarray14_uart3_rx_char_dupe2 = irqarray14_enable_storage[6];
assign irqarray14_uart3_err_dupe2 = irqarray14_enable_storage[7];
assign irqarray14_trng_done_dupe2 = irqarray14_enable_storage[8];
assign irqarray14_nc_b14s92 = irqarray14_enable_storage[9];
assign irqarray14_nc_b14s102 = irqarray14_enable_storage[10];
assign irqarray14_nc_b14s112 = irqarray14_enable_storage[11];
assign irqarray14_nc_b14s122 = irqarray14_enable_storage[12];
assign irqarray14_nc_b14s132 = irqarray14_enable_storage[13];
assign irqarray14_nc_b14s142 = irqarray14_enable_storage[14];
assign irqarray14_nc_b14s152 = irqarray14_enable_storage[15];
assign csrbank9_ev_enable0_w = irqarray14_enable_storage[15:0];
assign csrbank10_sel = (interface10_bank_bus_adr[15:10] == 4'd11);
assign csrbank10_re = interface10_bank_bus_re;
assign csrbank10_ev_soft0_r = interface10_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank10_ev_soft0_re <= 1'd0;
    csrbank10_ev_soft0_we <= 1'd0;
    if ((csrbank10_sel & (interface10_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank10_ev_soft0_re <= interface10_bank_bus_we;
        csrbank10_ev_soft0_we <= csrbank10_re;
    end
end
assign csrbank10_ev_edge_triggered0_r = interface10_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank10_ev_edge_triggered0_we <= 1'd0;
    csrbank10_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank10_sel & (interface10_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank10_ev_edge_triggered0_re <= interface10_bank_bus_we;
        csrbank10_ev_edge_triggered0_we <= csrbank10_re;
    end
end
assign csrbank10_ev_polarity0_r = interface10_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank10_ev_polarity0_we <= 1'd0;
    csrbank10_ev_polarity0_re <= 1'd0;
    if ((csrbank10_sel & (interface10_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank10_ev_polarity0_re <= interface10_bank_bus_we;
        csrbank10_ev_polarity0_we <= csrbank10_re;
    end
end
assign csrbank10_ev_status_r = interface10_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank10_ev_status_re <= 1'd0;
    csrbank10_ev_status_we <= 1'd0;
    if ((csrbank10_sel & (interface10_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank10_ev_status_re <= interface10_bank_bus_we;
        csrbank10_ev_status_we <= csrbank10_re;
    end
end
assign csrbank10_ev_pending_r = interface10_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank10_ev_pending_we <= 1'd0;
    csrbank10_ev_pending_re <= 1'd0;
    if ((csrbank10_sel & (interface10_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank10_ev_pending_re <= interface10_bank_bus_we;
        csrbank10_ev_pending_we <= csrbank10_re;
    end
end
assign csrbank10_ev_enable0_r = interface10_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank10_ev_enable0_we <= 1'd0;
    csrbank10_ev_enable0_re <= 1'd0;
    if ((csrbank10_sel & (interface10_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank10_ev_enable0_re <= interface10_bank_bus_we;
        csrbank10_ev_enable0_we <= csrbank10_re;
    end
end
always @(*) begin
    irqarray15_trigger <= 16'd0;
    if (irqarray15_soft_re) begin
        irqarray15_trigger <= irqarray15_soft_storage[15:0];
    end
end
assign csrbank10_ev_soft0_w = irqarray15_soft_storage[15:0];
assign irqarray15_use_edge = irqarray15_edge_triggered_storage[15:0];
assign csrbank10_ev_edge_triggered0_w = irqarray15_edge_triggered_storage[15:0];
assign irqarray15_rising = irqarray15_polarity_storage[15:0];
assign csrbank10_ev_polarity0_w = irqarray15_polarity_storage[15:0];
always @(*) begin
    irqarray15_status_status <= 16'd0;
    irqarray15_status_status[0] <= irqarray15_sec00;
    irqarray15_status_status[1] <= irqarray15_nc_b15s10;
    irqarray15_status_status[2] <= irqarray15_nc_b15s20;
    irqarray15_status_status[3] <= irqarray15_nc_b15s30;
    irqarray15_status_status[4] <= irqarray15_nc_b15s40;
    irqarray15_status_status[5] <= irqarray15_nc_b15s50;
    irqarray15_status_status[6] <= irqarray15_nc_b15s60;
    irqarray15_status_status[7] <= irqarray15_nc_b15s70;
    irqarray15_status_status[8] <= irqarray15_nc_b15s80;
    irqarray15_status_status[9] <= irqarray15_nc_b15s90;
    irqarray15_status_status[10] <= irqarray15_nc_b15s100;
    irqarray15_status_status[11] <= irqarray15_nc_b15s110;
    irqarray15_status_status[12] <= irqarray15_nc_b15s120;
    irqarray15_status_status[13] <= irqarray15_nc_b15s130;
    irqarray15_status_status[14] <= irqarray15_nc_b15s140;
    irqarray15_status_status[15] <= irqarray15_nc_b15s150;
end
assign csrbank10_ev_status_w = irqarray15_status_status[15:0];
assign irqarray15_status_we = csrbank10_ev_status_we;
always @(*) begin
    irqarray15_pending_status <= 16'd0;
    irqarray15_pending_status[0] <= irqarray15_sec01;
    irqarray15_pending_status[1] <= irqarray15_nc_b15s11;
    irqarray15_pending_status[2] <= irqarray15_nc_b15s21;
    irqarray15_pending_status[3] <= irqarray15_nc_b15s31;
    irqarray15_pending_status[4] <= irqarray15_nc_b15s41;
    irqarray15_pending_status[5] <= irqarray15_nc_b15s51;
    irqarray15_pending_status[6] <= irqarray15_nc_b15s61;
    irqarray15_pending_status[7] <= irqarray15_nc_b15s71;
    irqarray15_pending_status[8] <= irqarray15_nc_b15s81;
    irqarray15_pending_status[9] <= irqarray15_nc_b15s91;
    irqarray15_pending_status[10] <= irqarray15_nc_b15s101;
    irqarray15_pending_status[11] <= irqarray15_nc_b15s111;
    irqarray15_pending_status[12] <= irqarray15_nc_b15s121;
    irqarray15_pending_status[13] <= irqarray15_nc_b15s131;
    irqarray15_pending_status[14] <= irqarray15_nc_b15s141;
    irqarray15_pending_status[15] <= irqarray15_nc_b15s151;
end
assign csrbank10_ev_pending_w = irqarray15_pending_status[15:0];
assign irqarray15_pending_we = csrbank10_ev_pending_we;
assign irqarray15_sec02 = irqarray15_enable_storage[0];
assign irqarray15_nc_b15s12 = irqarray15_enable_storage[1];
assign irqarray15_nc_b15s22 = irqarray15_enable_storage[2];
assign irqarray15_nc_b15s32 = irqarray15_enable_storage[3];
assign irqarray15_nc_b15s42 = irqarray15_enable_storage[4];
assign irqarray15_nc_b15s52 = irqarray15_enable_storage[5];
assign irqarray15_nc_b15s62 = irqarray15_enable_storage[6];
assign irqarray15_nc_b15s72 = irqarray15_enable_storage[7];
assign irqarray15_nc_b15s82 = irqarray15_enable_storage[8];
assign irqarray15_nc_b15s92 = irqarray15_enable_storage[9];
assign irqarray15_nc_b15s102 = irqarray15_enable_storage[10];
assign irqarray15_nc_b15s112 = irqarray15_enable_storage[11];
assign irqarray15_nc_b15s122 = irqarray15_enable_storage[12];
assign irqarray15_nc_b15s132 = irqarray15_enable_storage[13];
assign irqarray15_nc_b15s142 = irqarray15_enable_storage[14];
assign irqarray15_nc_b15s152 = irqarray15_enable_storage[15];
assign csrbank10_ev_enable0_w = irqarray15_enable_storage[15:0];
assign csrbank11_sel = (interface11_bank_bus_adr[15:10] == 4'd12);
assign csrbank11_re = interface11_bank_bus_re;
assign csrbank11_ev_soft0_r = interface11_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank11_ev_soft0_re <= 1'd0;
    csrbank11_ev_soft0_we <= 1'd0;
    if ((csrbank11_sel & (interface11_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank11_ev_soft0_re <= interface11_bank_bus_we;
        csrbank11_ev_soft0_we <= csrbank11_re;
    end
end
assign csrbank11_ev_edge_triggered0_r = interface11_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank11_ev_edge_triggered0_we <= 1'd0;
    csrbank11_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank11_sel & (interface11_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank11_ev_edge_triggered0_re <= interface11_bank_bus_we;
        csrbank11_ev_edge_triggered0_we <= csrbank11_re;
    end
end
assign csrbank11_ev_polarity0_r = interface11_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank11_ev_polarity0_we <= 1'd0;
    csrbank11_ev_polarity0_re <= 1'd0;
    if ((csrbank11_sel & (interface11_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank11_ev_polarity0_re <= interface11_bank_bus_we;
        csrbank11_ev_polarity0_we <= csrbank11_re;
    end
end
assign csrbank11_ev_status_r = interface11_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank11_ev_status_re <= 1'd0;
    csrbank11_ev_status_we <= 1'd0;
    if ((csrbank11_sel & (interface11_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank11_ev_status_re <= interface11_bank_bus_we;
        csrbank11_ev_status_we <= csrbank11_re;
    end
end
assign csrbank11_ev_pending_r = interface11_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank11_ev_pending_we <= 1'd0;
    csrbank11_ev_pending_re <= 1'd0;
    if ((csrbank11_sel & (interface11_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank11_ev_pending_re <= interface11_bank_bus_we;
        csrbank11_ev_pending_we <= csrbank11_re;
    end
end
assign csrbank11_ev_enable0_r = interface11_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank11_ev_enable0_we <= 1'd0;
    csrbank11_ev_enable0_re <= 1'd0;
    if ((csrbank11_sel & (interface11_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank11_ev_enable0_re <= interface11_bank_bus_we;
        csrbank11_ev_enable0_we <= csrbank11_re;
    end
end
always @(*) begin
    irqarray16_trigger <= 16'd0;
    if (irqarray16_soft_re) begin
        irqarray16_trigger <= irqarray16_soft_storage[15:0];
    end
end
assign csrbank11_ev_soft0_w = irqarray16_soft_storage[15:0];
assign irqarray16_use_edge = irqarray16_edge_triggered_storage[15:0];
assign csrbank11_ev_edge_triggered0_w = irqarray16_edge_triggered_storage[15:0];
assign irqarray16_rising = irqarray16_polarity_storage[15:0];
assign csrbank11_ev_polarity0_w = irqarray16_polarity_storage[15:0];
always @(*) begin
    irqarray16_status_status <= 16'd0;
    irqarray16_status_status[0] <= irqarray16_cam_rx_dupe0;
    irqarray16_status_status[1] <= irqarray16_i2s_rx_dupe0;
    irqarray16_status_status[2] <= irqarray16_i2s_tx_dupe0;
    irqarray16_status_status[3] <= irqarray16_nc_b16s30;
    irqarray16_status_status[4] <= irqarray16_spim1_rx_dupe0;
    irqarray16_status_status[5] <= irqarray16_spim1_tx_dupe0;
    irqarray16_status_status[6] <= irqarray16_spim1_cmd_dupe0;
    irqarray16_status_status[7] <= irqarray16_spim1_eot_dupe0;
    irqarray16_status_status[8] <= irqarray16_spim2_rx_dupe0;
    irqarray16_status_status[9] <= irqarray16_spim2_tx_dupe0;
    irqarray16_status_status[10] <= irqarray16_spim2_cmd_dupe0;
    irqarray16_status_status[11] <= irqarray16_spim2_eot_dupe0;
    irqarray16_status_status[12] <= irqarray16_i2c0_rx_dupe0;
    irqarray16_status_status[13] <= irqarray16_i2c0_tx_dupe0;
    irqarray16_status_status[14] <= irqarray16_i2c0_cmd_dupe0;
    irqarray16_status_status[15] <= irqarray16_i2c0_eot_dupe0;
end
assign csrbank11_ev_status_w = irqarray16_status_status[15:0];
assign irqarray16_status_we = csrbank11_ev_status_we;
always @(*) begin
    irqarray16_pending_status <= 16'd0;
    irqarray16_pending_status[0] <= irqarray16_cam_rx_dupe1;
    irqarray16_pending_status[1] <= irqarray16_i2s_rx_dupe1;
    irqarray16_pending_status[2] <= irqarray16_i2s_tx_dupe1;
    irqarray16_pending_status[3] <= irqarray16_nc_b16s31;
    irqarray16_pending_status[4] <= irqarray16_spim1_rx_dupe1;
    irqarray16_pending_status[5] <= irqarray16_spim1_tx_dupe1;
    irqarray16_pending_status[6] <= irqarray16_spim1_cmd_dupe1;
    irqarray16_pending_status[7] <= irqarray16_spim1_eot_dupe1;
    irqarray16_pending_status[8] <= irqarray16_spim2_rx_dupe1;
    irqarray16_pending_status[9] <= irqarray16_spim2_tx_dupe1;
    irqarray16_pending_status[10] <= irqarray16_spim2_cmd_dupe1;
    irqarray16_pending_status[11] <= irqarray16_spim2_eot_dupe1;
    irqarray16_pending_status[12] <= irqarray16_i2c0_rx_dupe1;
    irqarray16_pending_status[13] <= irqarray16_i2c0_tx_dupe1;
    irqarray16_pending_status[14] <= irqarray16_i2c0_cmd_dupe1;
    irqarray16_pending_status[15] <= irqarray16_i2c0_eot_dupe1;
end
assign csrbank11_ev_pending_w = irqarray16_pending_status[15:0];
assign irqarray16_pending_we = csrbank11_ev_pending_we;
assign irqarray16_cam_rx_dupe2 = irqarray16_enable_storage[0];
assign irqarray16_i2s_rx_dupe2 = irqarray16_enable_storage[1];
assign irqarray16_i2s_tx_dupe2 = irqarray16_enable_storage[2];
assign irqarray16_nc_b16s32 = irqarray16_enable_storage[3];
assign irqarray16_spim1_rx_dupe2 = irqarray16_enable_storage[4];
assign irqarray16_spim1_tx_dupe2 = irqarray16_enable_storage[5];
assign irqarray16_spim1_cmd_dupe2 = irqarray16_enable_storage[6];
assign irqarray16_spim1_eot_dupe2 = irqarray16_enable_storage[7];
assign irqarray16_spim2_rx_dupe2 = irqarray16_enable_storage[8];
assign irqarray16_spim2_tx_dupe2 = irqarray16_enable_storage[9];
assign irqarray16_spim2_cmd_dupe2 = irqarray16_enable_storage[10];
assign irqarray16_spim2_eot_dupe2 = irqarray16_enable_storage[11];
assign irqarray16_i2c0_rx_dupe2 = irqarray16_enable_storage[12];
assign irqarray16_i2c0_tx_dupe2 = irqarray16_enable_storage[13];
assign irqarray16_i2c0_cmd_dupe2 = irqarray16_enable_storage[14];
assign irqarray16_i2c0_eot_dupe2 = irqarray16_enable_storage[15];
assign csrbank11_ev_enable0_w = irqarray16_enable_storage[15:0];
assign csrbank12_sel = (interface12_bank_bus_adr[15:10] == 4'd13);
assign csrbank12_re = interface12_bank_bus_re;
assign csrbank12_ev_soft0_r = interface12_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank12_ev_soft0_re <= 1'd0;
    csrbank12_ev_soft0_we <= 1'd0;
    if ((csrbank12_sel & (interface12_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank12_ev_soft0_re <= interface12_bank_bus_we;
        csrbank12_ev_soft0_we <= csrbank12_re;
    end
end
assign csrbank12_ev_edge_triggered0_r = interface12_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank12_ev_edge_triggered0_we <= 1'd0;
    csrbank12_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank12_sel & (interface12_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank12_ev_edge_triggered0_re <= interface12_bank_bus_we;
        csrbank12_ev_edge_triggered0_we <= csrbank12_re;
    end
end
assign csrbank12_ev_polarity0_r = interface12_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank12_ev_polarity0_we <= 1'd0;
    csrbank12_ev_polarity0_re <= 1'd0;
    if ((csrbank12_sel & (interface12_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank12_ev_polarity0_re <= interface12_bank_bus_we;
        csrbank12_ev_polarity0_we <= csrbank12_re;
    end
end
assign csrbank12_ev_status_r = interface12_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank12_ev_status_re <= 1'd0;
    csrbank12_ev_status_we <= 1'd0;
    if ((csrbank12_sel & (interface12_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank12_ev_status_re <= interface12_bank_bus_we;
        csrbank12_ev_status_we <= csrbank12_re;
    end
end
assign csrbank12_ev_pending_r = interface12_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank12_ev_pending_we <= 1'd0;
    csrbank12_ev_pending_re <= 1'd0;
    if ((csrbank12_sel & (interface12_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank12_ev_pending_re <= interface12_bank_bus_we;
        csrbank12_ev_pending_we <= csrbank12_re;
    end
end
assign csrbank12_ev_enable0_r = interface12_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank12_ev_enable0_we <= 1'd0;
    csrbank12_ev_enable0_re <= 1'd0;
    if ((csrbank12_sel & (interface12_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank12_ev_enable0_re <= interface12_bank_bus_we;
        csrbank12_ev_enable0_we <= csrbank12_re;
    end
end
always @(*) begin
    irqarray17_trigger <= 16'd0;
    if (irqarray17_soft_re) begin
        irqarray17_trigger <= irqarray17_soft_storage[15:0];
    end
end
assign csrbank12_ev_soft0_w = irqarray17_soft_storage[15:0];
assign irqarray17_use_edge = irqarray17_edge_triggered_storage[15:0];
assign csrbank12_ev_edge_triggered0_w = irqarray17_edge_triggered_storage[15:0];
assign irqarray17_rising = irqarray17_polarity_storage[15:0];
assign csrbank12_ev_polarity0_w = irqarray17_polarity_storage[15:0];
always @(*) begin
    irqarray17_status_status <= 16'd0;
    irqarray17_status_status[0] <= irqarray17_i2c1_rx_dupe0;
    irqarray17_status_status[1] <= irqarray17_i2c1_tx_dupe0;
    irqarray17_status_status[2] <= irqarray17_i2c1_cmd_dupe0;
    irqarray17_status_status[3] <= irqarray17_i2c1_eot_dupe0;
    irqarray17_status_status[4] <= irqarray17_pioirq0_dupe0;
    irqarray17_status_status[5] <= irqarray17_pioirq1_dupe0;
    irqarray17_status_status[6] <= irqarray17_pioirq2_dupe0;
    irqarray17_status_status[7] <= irqarray17_pioirq3_dupe0;
    irqarray17_status_status[8] <= irqarray17_qfcirq_dupe0;
    irqarray17_status_status[9] <= irqarray17_adc_rx_dupe0;
    irqarray17_status_status[10] <= irqarray17_ioxirq_dupe0;
    irqarray17_status_status[11] <= irqarray17_sddcirq_dupe0;
    irqarray17_status_status[12] <= irqarray17_nc_b17s120;
    irqarray17_status_status[13] <= irqarray17_nc_b17s130;
    irqarray17_status_status[14] <= irqarray17_nc_b17s140;
    irqarray17_status_status[15] <= irqarray17_nc_b17s150;
end
assign csrbank12_ev_status_w = irqarray17_status_status[15:0];
assign irqarray17_status_we = csrbank12_ev_status_we;
always @(*) begin
    irqarray17_pending_status <= 16'd0;
    irqarray17_pending_status[0] <= irqarray17_i2c1_rx_dupe1;
    irqarray17_pending_status[1] <= irqarray17_i2c1_tx_dupe1;
    irqarray17_pending_status[2] <= irqarray17_i2c1_cmd_dupe1;
    irqarray17_pending_status[3] <= irqarray17_i2c1_eot_dupe1;
    irqarray17_pending_status[4] <= irqarray17_pioirq0_dupe1;
    irqarray17_pending_status[5] <= irqarray17_pioirq1_dupe1;
    irqarray17_pending_status[6] <= irqarray17_pioirq2_dupe1;
    irqarray17_pending_status[7] <= irqarray17_pioirq3_dupe1;
    irqarray17_pending_status[8] <= irqarray17_qfcirq_dupe1;
    irqarray17_pending_status[9] <= irqarray17_adc_rx_dupe1;
    irqarray17_pending_status[10] <= irqarray17_ioxirq_dupe1;
    irqarray17_pending_status[11] <= irqarray17_sddcirq_dupe1;
    irqarray17_pending_status[12] <= irqarray17_nc_b17s121;
    irqarray17_pending_status[13] <= irqarray17_nc_b17s131;
    irqarray17_pending_status[14] <= irqarray17_nc_b17s141;
    irqarray17_pending_status[15] <= irqarray17_nc_b17s151;
end
assign csrbank12_ev_pending_w = irqarray17_pending_status[15:0];
assign irqarray17_pending_we = csrbank12_ev_pending_we;
assign irqarray17_i2c1_rx_dupe2 = irqarray17_enable_storage[0];
assign irqarray17_i2c1_tx_dupe2 = irqarray17_enable_storage[1];
assign irqarray17_i2c1_cmd_dupe2 = irqarray17_enable_storage[2];
assign irqarray17_i2c1_eot_dupe2 = irqarray17_enable_storage[3];
assign irqarray17_pioirq0_dupe2 = irqarray17_enable_storage[4];
assign irqarray17_pioirq1_dupe2 = irqarray17_enable_storage[5];
assign irqarray17_pioirq2_dupe2 = irqarray17_enable_storage[6];
assign irqarray17_pioirq3_dupe2 = irqarray17_enable_storage[7];
assign irqarray17_qfcirq_dupe2 = irqarray17_enable_storage[8];
assign irqarray17_adc_rx_dupe2 = irqarray17_enable_storage[9];
assign irqarray17_ioxirq_dupe2 = irqarray17_enable_storage[10];
assign irqarray17_sddcirq_dupe2 = irqarray17_enable_storage[11];
assign irqarray17_nc_b17s122 = irqarray17_enable_storage[12];
assign irqarray17_nc_b17s132 = irqarray17_enable_storage[13];
assign irqarray17_nc_b17s142 = irqarray17_enable_storage[14];
assign irqarray17_nc_b17s152 = irqarray17_enable_storage[15];
assign csrbank12_ev_enable0_w = irqarray17_enable_storage[15:0];
assign csrbank13_sel = (interface13_bank_bus_adr[15:10] == 4'd14);
assign csrbank13_re = interface13_bank_bus_re;
assign csrbank13_ev_soft0_r = interface13_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank13_ev_soft0_re <= 1'd0;
    csrbank13_ev_soft0_we <= 1'd0;
    if ((csrbank13_sel & (interface13_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank13_ev_soft0_re <= interface13_bank_bus_we;
        csrbank13_ev_soft0_we <= csrbank13_re;
    end
end
assign csrbank13_ev_edge_triggered0_r = interface13_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank13_ev_edge_triggered0_we <= 1'd0;
    csrbank13_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank13_sel & (interface13_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank13_ev_edge_triggered0_re <= interface13_bank_bus_we;
        csrbank13_ev_edge_triggered0_we <= csrbank13_re;
    end
end
assign csrbank13_ev_polarity0_r = interface13_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank13_ev_polarity0_we <= 1'd0;
    csrbank13_ev_polarity0_re <= 1'd0;
    if ((csrbank13_sel & (interface13_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank13_ev_polarity0_re <= interface13_bank_bus_we;
        csrbank13_ev_polarity0_we <= csrbank13_re;
    end
end
assign csrbank13_ev_status_r = interface13_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank13_ev_status_re <= 1'd0;
    csrbank13_ev_status_we <= 1'd0;
    if ((csrbank13_sel & (interface13_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank13_ev_status_re <= interface13_bank_bus_we;
        csrbank13_ev_status_we <= csrbank13_re;
    end
end
assign csrbank13_ev_pending_r = interface13_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank13_ev_pending_we <= 1'd0;
    csrbank13_ev_pending_re <= 1'd0;
    if ((csrbank13_sel & (interface13_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank13_ev_pending_re <= interface13_bank_bus_we;
        csrbank13_ev_pending_we <= csrbank13_re;
    end
end
assign csrbank13_ev_enable0_r = interface13_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank13_ev_enable0_we <= 1'd0;
    csrbank13_ev_enable0_re <= 1'd0;
    if ((csrbank13_sel & (interface13_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank13_ev_enable0_re <= interface13_bank_bus_we;
        csrbank13_ev_enable0_we <= csrbank13_re;
    end
end
always @(*) begin
    irqarray18_trigger <= 16'd0;
    if (irqarray18_soft_re) begin
        irqarray18_trigger <= irqarray18_soft_storage[15:0];
    end
end
assign csrbank13_ev_soft0_w = irqarray18_soft_storage[15:0];
assign irqarray18_use_edge = irqarray18_edge_triggered_storage[15:0];
assign csrbank13_ev_edge_triggered0_w = irqarray18_edge_triggered_storage[15:0];
assign irqarray18_rising = irqarray18_polarity_storage[15:0];
assign csrbank13_ev_polarity0_w = irqarray18_polarity_storage[15:0];
always @(*) begin
    irqarray18_status_status <= 16'd0;
    irqarray18_status_status[0] <= irqarray18_pioirq0_dupe0;
    irqarray18_status_status[1] <= irqarray18_pioirq1_dupe0;
    irqarray18_status_status[2] <= irqarray18_pioirq2_dupe0;
    irqarray18_status_status[3] <= irqarray18_pioirq3_dupe0;
    irqarray18_status_status[4] <= irqarray18_i2c2_rx_dupe0;
    irqarray18_status_status[5] <= irqarray18_i2c2_tx_dupe0;
    irqarray18_status_status[6] <= irqarray18_i2c2_cmd_dupe0;
    irqarray18_status_status[7] <= irqarray18_i2c2_eot_dupe0;
    irqarray18_status_status[8] <= irqarray18_i2c0_nack_dupe0;
    irqarray18_status_status[9] <= irqarray18_i2c1_nack_dupe0;
    irqarray18_status_status[10] <= irqarray18_i2c2_nack_dupe0;
    irqarray18_status_status[11] <= irqarray18_i2c0_err_dupe0;
    irqarray18_status_status[12] <= irqarray18_i2c1_err_dupe0;
    irqarray18_status_status[13] <= irqarray18_i2c2_err_dupe0;
    irqarray18_status_status[14] <= irqarray18_ioxirq_dupe0;
    irqarray18_status_status[15] <= irqarray18_cam_rx_dupe0;
end
assign csrbank13_ev_status_w = irqarray18_status_status[15:0];
assign irqarray18_status_we = csrbank13_ev_status_we;
always @(*) begin
    irqarray18_pending_status <= 16'd0;
    irqarray18_pending_status[0] <= irqarray18_pioirq0_dupe1;
    irqarray18_pending_status[1] <= irqarray18_pioirq1_dupe1;
    irqarray18_pending_status[2] <= irqarray18_pioirq2_dupe1;
    irqarray18_pending_status[3] <= irqarray18_pioirq3_dupe1;
    irqarray18_pending_status[4] <= irqarray18_i2c2_rx_dupe1;
    irqarray18_pending_status[5] <= irqarray18_i2c2_tx_dupe1;
    irqarray18_pending_status[6] <= irqarray18_i2c2_cmd_dupe1;
    irqarray18_pending_status[7] <= irqarray18_i2c2_eot_dupe1;
    irqarray18_pending_status[8] <= irqarray18_i2c0_nack_dupe1;
    irqarray18_pending_status[9] <= irqarray18_i2c1_nack_dupe1;
    irqarray18_pending_status[10] <= irqarray18_i2c2_nack_dupe1;
    irqarray18_pending_status[11] <= irqarray18_i2c0_err_dupe1;
    irqarray18_pending_status[12] <= irqarray18_i2c1_err_dupe1;
    irqarray18_pending_status[13] <= irqarray18_i2c2_err_dupe1;
    irqarray18_pending_status[14] <= irqarray18_ioxirq_dupe1;
    irqarray18_pending_status[15] <= irqarray18_cam_rx_dupe1;
end
assign csrbank13_ev_pending_w = irqarray18_pending_status[15:0];
assign irqarray18_pending_we = csrbank13_ev_pending_we;
assign irqarray18_pioirq0_dupe2 = irqarray18_enable_storage[0];
assign irqarray18_pioirq1_dupe2 = irqarray18_enable_storage[1];
assign irqarray18_pioirq2_dupe2 = irqarray18_enable_storage[2];
assign irqarray18_pioirq3_dupe2 = irqarray18_enable_storage[3];
assign irqarray18_i2c2_rx_dupe2 = irqarray18_enable_storage[4];
assign irqarray18_i2c2_tx_dupe2 = irqarray18_enable_storage[5];
assign irqarray18_i2c2_cmd_dupe2 = irqarray18_enable_storage[6];
assign irqarray18_i2c2_eot_dupe2 = irqarray18_enable_storage[7];
assign irqarray18_i2c0_nack_dupe2 = irqarray18_enable_storage[8];
assign irqarray18_i2c1_nack_dupe2 = irqarray18_enable_storage[9];
assign irqarray18_i2c2_nack_dupe2 = irqarray18_enable_storage[10];
assign irqarray18_i2c0_err_dupe2 = irqarray18_enable_storage[11];
assign irqarray18_i2c1_err_dupe2 = irqarray18_enable_storage[12];
assign irqarray18_i2c2_err_dupe2 = irqarray18_enable_storage[13];
assign irqarray18_ioxirq_dupe2 = irqarray18_enable_storage[14];
assign irqarray18_cam_rx_dupe2 = irqarray18_enable_storage[15];
assign csrbank13_ev_enable0_w = irqarray18_enable_storage[15:0];
assign csrbank14_sel = (interface14_bank_bus_adr[15:10] == 4'd15);
assign csrbank14_re = interface14_bank_bus_re;
assign csrbank14_ev_soft0_r = interface14_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank14_ev_soft0_re <= 1'd0;
    csrbank14_ev_soft0_we <= 1'd0;
    if ((csrbank14_sel & (interface14_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank14_ev_soft0_re <= interface14_bank_bus_we;
        csrbank14_ev_soft0_we <= csrbank14_re;
    end
end
assign csrbank14_ev_edge_triggered0_r = interface14_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank14_ev_edge_triggered0_we <= 1'd0;
    csrbank14_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank14_sel & (interface14_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank14_ev_edge_triggered0_re <= interface14_bank_bus_we;
        csrbank14_ev_edge_triggered0_we <= csrbank14_re;
    end
end
assign csrbank14_ev_polarity0_r = interface14_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank14_ev_polarity0_we <= 1'd0;
    csrbank14_ev_polarity0_re <= 1'd0;
    if ((csrbank14_sel & (interface14_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank14_ev_polarity0_re <= interface14_bank_bus_we;
        csrbank14_ev_polarity0_we <= csrbank14_re;
    end
end
assign csrbank14_ev_status_r = interface14_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank14_ev_status_re <= 1'd0;
    csrbank14_ev_status_we <= 1'd0;
    if ((csrbank14_sel & (interface14_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank14_ev_status_re <= interface14_bank_bus_we;
        csrbank14_ev_status_we <= csrbank14_re;
    end
end
assign csrbank14_ev_pending_r = interface14_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank14_ev_pending_we <= 1'd0;
    csrbank14_ev_pending_re <= 1'd0;
    if ((csrbank14_sel & (interface14_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank14_ev_pending_re <= interface14_bank_bus_we;
        csrbank14_ev_pending_we <= csrbank14_re;
    end
end
assign csrbank14_ev_enable0_r = interface14_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank14_ev_enable0_we <= 1'd0;
    csrbank14_ev_enable0_re <= 1'd0;
    if ((csrbank14_sel & (interface14_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank14_ev_enable0_re <= interface14_bank_bus_we;
        csrbank14_ev_enable0_we <= csrbank14_re;
    end
end
always @(*) begin
    irqarray19_trigger <= 16'd0;
    if (irqarray19_soft_re) begin
        irqarray19_trigger <= irqarray19_soft_storage[15:0];
    end
end
assign csrbank14_ev_soft0_w = irqarray19_soft_storage[15:0];
assign irqarray19_use_edge = irqarray19_edge_triggered_storage[15:0];
assign csrbank14_ev_edge_triggered0_w = irqarray19_edge_triggered_storage[15:0];
assign irqarray19_rising = irqarray19_polarity_storage[15:0];
assign csrbank14_ev_polarity0_w = irqarray19_polarity_storage[15:0];
always @(*) begin
    irqarray19_status_status <= 16'd0;
    irqarray19_status_status[0] <= irqarray19_mbox_irq_available_dupe0;
    irqarray19_status_status[1] <= irqarray19_mbox_irq_abort_init_dupe0;
    irqarray19_status_status[2] <= irqarray19_mbox_irq_done_dupe0;
    irqarray19_status_status[3] <= irqarray19_mbox_irq_error_dupe0;
    irqarray19_status_status[4] <= irqarray19_pioirq0_dupe0;
    irqarray19_status_status[5] <= irqarray19_pioirq1_dupe0;
    irqarray19_status_status[6] <= irqarray19_pioirq2_dupe0;
    irqarray19_status_status[7] <= irqarray19_pioirq3_dupe0;
    irqarray19_status_status[8] <= irqarray19_sdio_rx_dupe0;
    irqarray19_status_status[9] <= irqarray19_sdio_tx_dupe0;
    irqarray19_status_status[10] <= irqarray19_sdio_eot_dupe0;
    irqarray19_status_status[11] <= irqarray19_sdio_err_dupe0;
    irqarray19_status_status[12] <= irqarray19_nc_b19s120;
    irqarray19_status_status[13] <= irqarray19_nc_b19s130;
    irqarray19_status_status[14] <= irqarray19_nc_b19s140;
    irqarray19_status_status[15] <= irqarray19_nc_b19s150;
end
assign csrbank14_ev_status_w = irqarray19_status_status[15:0];
assign irqarray19_status_we = csrbank14_ev_status_we;
always @(*) begin
    irqarray19_pending_status <= 16'd0;
    irqarray19_pending_status[0] <= irqarray19_mbox_irq_available_dupe1;
    irqarray19_pending_status[1] <= irqarray19_mbox_irq_abort_init_dupe1;
    irqarray19_pending_status[2] <= irqarray19_mbox_irq_done_dupe1;
    irqarray19_pending_status[3] <= irqarray19_mbox_irq_error_dupe1;
    irqarray19_pending_status[4] <= irqarray19_pioirq0_dupe1;
    irqarray19_pending_status[5] <= irqarray19_pioirq1_dupe1;
    irqarray19_pending_status[6] <= irqarray19_pioirq2_dupe1;
    irqarray19_pending_status[7] <= irqarray19_pioirq3_dupe1;
    irqarray19_pending_status[8] <= irqarray19_sdio_rx_dupe1;
    irqarray19_pending_status[9] <= irqarray19_sdio_tx_dupe1;
    irqarray19_pending_status[10] <= irqarray19_sdio_eot_dupe1;
    irqarray19_pending_status[11] <= irqarray19_sdio_err_dupe1;
    irqarray19_pending_status[12] <= irqarray19_nc_b19s121;
    irqarray19_pending_status[13] <= irqarray19_nc_b19s131;
    irqarray19_pending_status[14] <= irqarray19_nc_b19s141;
    irqarray19_pending_status[15] <= irqarray19_nc_b19s151;
end
assign csrbank14_ev_pending_w = irqarray19_pending_status[15:0];
assign irqarray19_pending_we = csrbank14_ev_pending_we;
assign irqarray19_mbox_irq_available_dupe2 = irqarray19_enable_storage[0];
assign irqarray19_mbox_irq_abort_init_dupe2 = irqarray19_enable_storage[1];
assign irqarray19_mbox_irq_done_dupe2 = irqarray19_enable_storage[2];
assign irqarray19_mbox_irq_error_dupe2 = irqarray19_enable_storage[3];
assign irqarray19_pioirq0_dupe2 = irqarray19_enable_storage[4];
assign irqarray19_pioirq1_dupe2 = irqarray19_enable_storage[5];
assign irqarray19_pioirq2_dupe2 = irqarray19_enable_storage[6];
assign irqarray19_pioirq3_dupe2 = irqarray19_enable_storage[7];
assign irqarray19_sdio_rx_dupe2 = irqarray19_enable_storage[8];
assign irqarray19_sdio_tx_dupe2 = irqarray19_enable_storage[9];
assign irqarray19_sdio_eot_dupe2 = irqarray19_enable_storage[10];
assign irqarray19_sdio_err_dupe2 = irqarray19_enable_storage[11];
assign irqarray19_nc_b19s122 = irqarray19_enable_storage[12];
assign irqarray19_nc_b19s132 = irqarray19_enable_storage[13];
assign irqarray19_nc_b19s142 = irqarray19_enable_storage[14];
assign irqarray19_nc_b19s152 = irqarray19_enable_storage[15];
assign csrbank14_ev_enable0_w = irqarray19_enable_storage[15:0];
assign csrbank15_sel = (interface15_bank_bus_adr[15:10] == 5'd16);
assign csrbank15_re = interface15_bank_bus_re;
assign csrbank15_ev_soft0_r = interface15_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank15_ev_soft0_re <= 1'd0;
    csrbank15_ev_soft0_we <= 1'd0;
    if ((csrbank15_sel & (interface15_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank15_ev_soft0_re <= interface15_bank_bus_we;
        csrbank15_ev_soft0_we <= csrbank15_re;
    end
end
assign csrbank15_ev_edge_triggered0_r = interface15_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank15_ev_edge_triggered0_we <= 1'd0;
    csrbank15_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank15_sel & (interface15_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank15_ev_edge_triggered0_re <= interface15_bank_bus_we;
        csrbank15_ev_edge_triggered0_we <= csrbank15_re;
    end
end
assign csrbank15_ev_polarity0_r = interface15_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank15_ev_polarity0_we <= 1'd0;
    csrbank15_ev_polarity0_re <= 1'd0;
    if ((csrbank15_sel & (interface15_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank15_ev_polarity0_re <= interface15_bank_bus_we;
        csrbank15_ev_polarity0_we <= csrbank15_re;
    end
end
assign csrbank15_ev_status_r = interface15_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank15_ev_status_re <= 1'd0;
    csrbank15_ev_status_we <= 1'd0;
    if ((csrbank15_sel & (interface15_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank15_ev_status_re <= interface15_bank_bus_we;
        csrbank15_ev_status_we <= csrbank15_re;
    end
end
assign csrbank15_ev_pending_r = interface15_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank15_ev_pending_we <= 1'd0;
    csrbank15_ev_pending_re <= 1'd0;
    if ((csrbank15_sel & (interface15_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank15_ev_pending_re <= interface15_bank_bus_we;
        csrbank15_ev_pending_we <= csrbank15_re;
    end
end
assign csrbank15_ev_enable0_r = interface15_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank15_ev_enable0_we <= 1'd0;
    csrbank15_ev_enable0_re <= 1'd0;
    if ((csrbank15_sel & (interface15_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank15_ev_enable0_re <= interface15_bank_bus_we;
        csrbank15_ev_enable0_we <= csrbank15_re;
    end
end
always @(*) begin
    irqarray2_trigger <= 16'd0;
    if (irqarray2_soft_re) begin
        irqarray2_trigger <= irqarray2_soft_storage[15:0];
    end
end
assign csrbank15_ev_soft0_w = irqarray2_soft_storage[15:0];
assign irqarray2_use_edge = irqarray2_edge_triggered_storage[15:0];
assign csrbank15_ev_edge_triggered0_w = irqarray2_edge_triggered_storage[15:0];
assign irqarray2_rising = irqarray2_polarity_storage[15:0];
assign csrbank15_ev_polarity0_w = irqarray2_polarity_storage[15:0];
always @(*) begin
    irqarray2_status_status <= 16'd0;
    irqarray2_status_status[0] <= irqarray2_qfcirq0;
    irqarray2_status_status[1] <= irqarray2_mdmairq0;
    irqarray2_status_status[2] <= irqarray2_mbox_irq_available0;
    irqarray2_status_status[3] <= irqarray2_mbox_irq_abort_init0;
    irqarray2_status_status[4] <= irqarray2_mbox_irq_done0;
    irqarray2_status_status[5] <= irqarray2_mbox_irq_error0;
    irqarray2_status_status[6] <= irqarray2_nc_b2s60;
    irqarray2_status_status[7] <= irqarray2_nc_b2s70;
    irqarray2_status_status[8] <= irqarray2_nc_b2s80;
    irqarray2_status_status[9] <= irqarray2_nc_b2s90;
    irqarray2_status_status[10] <= irqarray2_nc_b2s100;
    irqarray2_status_status[11] <= irqarray2_nc_b2s110;
    irqarray2_status_status[12] <= irqarray2_nc_b2s120;
    irqarray2_status_status[13] <= irqarray2_nc_b2s130;
    irqarray2_status_status[14] <= irqarray2_nc_b2s140;
    irqarray2_status_status[15] <= irqarray2_aowkupint0;
end
assign csrbank15_ev_status_w = irqarray2_status_status[15:0];
assign irqarray2_status_we = csrbank15_ev_status_we;
always @(*) begin
    irqarray2_pending_status <= 16'd0;
    irqarray2_pending_status[0] <= irqarray2_qfcirq1;
    irqarray2_pending_status[1] <= irqarray2_mdmairq1;
    irqarray2_pending_status[2] <= irqarray2_mbox_irq_available1;
    irqarray2_pending_status[3] <= irqarray2_mbox_irq_abort_init1;
    irqarray2_pending_status[4] <= irqarray2_mbox_irq_done1;
    irqarray2_pending_status[5] <= irqarray2_mbox_irq_error1;
    irqarray2_pending_status[6] <= irqarray2_nc_b2s61;
    irqarray2_pending_status[7] <= irqarray2_nc_b2s71;
    irqarray2_pending_status[8] <= irqarray2_nc_b2s81;
    irqarray2_pending_status[9] <= irqarray2_nc_b2s91;
    irqarray2_pending_status[10] <= irqarray2_nc_b2s101;
    irqarray2_pending_status[11] <= irqarray2_nc_b2s111;
    irqarray2_pending_status[12] <= irqarray2_nc_b2s121;
    irqarray2_pending_status[13] <= irqarray2_nc_b2s131;
    irqarray2_pending_status[14] <= irqarray2_nc_b2s141;
    irqarray2_pending_status[15] <= irqarray2_aowkupint1;
end
assign csrbank15_ev_pending_w = irqarray2_pending_status[15:0];
assign irqarray2_pending_we = csrbank15_ev_pending_we;
assign irqarray2_qfcirq2 = irqarray2_enable_storage[0];
assign irqarray2_mdmairq2 = irqarray2_enable_storage[1];
assign irqarray2_mbox_irq_available2 = irqarray2_enable_storage[2];
assign irqarray2_mbox_irq_abort_init2 = irqarray2_enable_storage[3];
assign irqarray2_mbox_irq_done2 = irqarray2_enable_storage[4];
assign irqarray2_mbox_irq_error2 = irqarray2_enable_storage[5];
assign irqarray2_nc_b2s62 = irqarray2_enable_storage[6];
assign irqarray2_nc_b2s72 = irqarray2_enable_storage[7];
assign irqarray2_nc_b2s82 = irqarray2_enable_storage[8];
assign irqarray2_nc_b2s92 = irqarray2_enable_storage[9];
assign irqarray2_nc_b2s102 = irqarray2_enable_storage[10];
assign irqarray2_nc_b2s112 = irqarray2_enable_storage[11];
assign irqarray2_nc_b2s122 = irqarray2_enable_storage[12];
assign irqarray2_nc_b2s132 = irqarray2_enable_storage[13];
assign irqarray2_nc_b2s142 = irqarray2_enable_storage[14];
assign irqarray2_aowkupint2 = irqarray2_enable_storage[15];
assign csrbank15_ev_enable0_w = irqarray2_enable_storage[15:0];
assign csrbank16_sel = (interface16_bank_bus_adr[15:10] == 5'd17);
assign csrbank16_re = interface16_bank_bus_re;
assign csrbank16_ev_soft0_r = interface16_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank16_ev_soft0_re <= 1'd0;
    csrbank16_ev_soft0_we <= 1'd0;
    if ((csrbank16_sel & (interface16_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank16_ev_soft0_re <= interface16_bank_bus_we;
        csrbank16_ev_soft0_we <= csrbank16_re;
    end
end
assign csrbank16_ev_edge_triggered0_r = interface16_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank16_ev_edge_triggered0_we <= 1'd0;
    csrbank16_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank16_sel & (interface16_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank16_ev_edge_triggered0_re <= interface16_bank_bus_we;
        csrbank16_ev_edge_triggered0_we <= csrbank16_re;
    end
end
assign csrbank16_ev_polarity0_r = interface16_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank16_ev_polarity0_we <= 1'd0;
    csrbank16_ev_polarity0_re <= 1'd0;
    if ((csrbank16_sel & (interface16_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank16_ev_polarity0_re <= interface16_bank_bus_we;
        csrbank16_ev_polarity0_we <= csrbank16_re;
    end
end
assign csrbank16_ev_status_r = interface16_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank16_ev_status_re <= 1'd0;
    csrbank16_ev_status_we <= 1'd0;
    if ((csrbank16_sel & (interface16_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank16_ev_status_re <= interface16_bank_bus_we;
        csrbank16_ev_status_we <= csrbank16_re;
    end
end
assign csrbank16_ev_pending_r = interface16_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank16_ev_pending_we <= 1'd0;
    csrbank16_ev_pending_re <= 1'd0;
    if ((csrbank16_sel & (interface16_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank16_ev_pending_re <= interface16_bank_bus_we;
        csrbank16_ev_pending_we <= csrbank16_re;
    end
end
assign csrbank16_ev_enable0_r = interface16_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank16_ev_enable0_we <= 1'd0;
    csrbank16_ev_enable0_re <= 1'd0;
    if ((csrbank16_sel & (interface16_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank16_ev_enable0_re <= interface16_bank_bus_we;
        csrbank16_ev_enable0_we <= csrbank16_re;
    end
end
always @(*) begin
    irqarray3_trigger <= 16'd0;
    if (irqarray3_soft_re) begin
        irqarray3_trigger <= irqarray3_soft_storage[15:0];
    end
end
assign csrbank16_ev_soft0_w = irqarray3_soft_storage[15:0];
assign irqarray3_use_edge = irqarray3_edge_triggered_storage[15:0];
assign csrbank16_ev_edge_triggered0_w = irqarray3_edge_triggered_storage[15:0];
assign irqarray3_rising = irqarray3_polarity_storage[15:0];
assign csrbank16_ev_polarity0_w = irqarray3_polarity_storage[15:0];
always @(*) begin
    irqarray3_status_status <= 16'd0;
    irqarray3_status_status[0] <= irqarray3_trng_done0;
    irqarray3_status_status[1] <= irqarray3_aes_done0;
    irqarray3_status_status[2] <= irqarray3_pke_done0;
    irqarray3_status_status[3] <= irqarray3_hash_done0;
    irqarray3_status_status[4] <= irqarray3_alu_done0;
    irqarray3_status_status[5] <= irqarray3_sdma_ichdone0;
    irqarray3_status_status[6] <= irqarray3_sdma_schdone0;
    irqarray3_status_status[7] <= irqarray3_sdma_xchdone0;
    irqarray3_status_status[8] <= irqarray3_nc_b3s80;
    irqarray3_status_status[9] <= irqarray3_nc_b3s90;
    irqarray3_status_status[10] <= irqarray3_nc_b3s100;
    irqarray3_status_status[11] <= irqarray3_nc_b3s110;
    irqarray3_status_status[12] <= irqarray3_nc_b3s120;
    irqarray3_status_status[13] <= irqarray3_nc_b3s130;
    irqarray3_status_status[14] <= irqarray3_nc_b3s140;
    irqarray3_status_status[15] <= irqarray3_nc_b3s150;
end
assign csrbank16_ev_status_w = irqarray3_status_status[15:0];
assign irqarray3_status_we = csrbank16_ev_status_we;
always @(*) begin
    irqarray3_pending_status <= 16'd0;
    irqarray3_pending_status[0] <= irqarray3_trng_done1;
    irqarray3_pending_status[1] <= irqarray3_aes_done1;
    irqarray3_pending_status[2] <= irqarray3_pke_done1;
    irqarray3_pending_status[3] <= irqarray3_hash_done1;
    irqarray3_pending_status[4] <= irqarray3_alu_done1;
    irqarray3_pending_status[5] <= irqarray3_sdma_ichdone1;
    irqarray3_pending_status[6] <= irqarray3_sdma_schdone1;
    irqarray3_pending_status[7] <= irqarray3_sdma_xchdone1;
    irqarray3_pending_status[8] <= irqarray3_nc_b3s81;
    irqarray3_pending_status[9] <= irqarray3_nc_b3s91;
    irqarray3_pending_status[10] <= irqarray3_nc_b3s101;
    irqarray3_pending_status[11] <= irqarray3_nc_b3s111;
    irqarray3_pending_status[12] <= irqarray3_nc_b3s121;
    irqarray3_pending_status[13] <= irqarray3_nc_b3s131;
    irqarray3_pending_status[14] <= irqarray3_nc_b3s141;
    irqarray3_pending_status[15] <= irqarray3_nc_b3s151;
end
assign csrbank16_ev_pending_w = irqarray3_pending_status[15:0];
assign irqarray3_pending_we = csrbank16_ev_pending_we;
assign irqarray3_trng_done2 = irqarray3_enable_storage[0];
assign irqarray3_aes_done2 = irqarray3_enable_storage[1];
assign irqarray3_pke_done2 = irqarray3_enable_storage[2];
assign irqarray3_hash_done2 = irqarray3_enable_storage[3];
assign irqarray3_alu_done2 = irqarray3_enable_storage[4];
assign irqarray3_sdma_ichdone2 = irqarray3_enable_storage[5];
assign irqarray3_sdma_schdone2 = irqarray3_enable_storage[6];
assign irqarray3_sdma_xchdone2 = irqarray3_enable_storage[7];
assign irqarray3_nc_b3s82 = irqarray3_enable_storage[8];
assign irqarray3_nc_b3s92 = irqarray3_enable_storage[9];
assign irqarray3_nc_b3s102 = irqarray3_enable_storage[10];
assign irqarray3_nc_b3s112 = irqarray3_enable_storage[11];
assign irqarray3_nc_b3s122 = irqarray3_enable_storage[12];
assign irqarray3_nc_b3s132 = irqarray3_enable_storage[13];
assign irqarray3_nc_b3s142 = irqarray3_enable_storage[14];
assign irqarray3_nc_b3s152 = irqarray3_enable_storage[15];
assign csrbank16_ev_enable0_w = irqarray3_enable_storage[15:0];
assign csrbank17_sel = (interface17_bank_bus_adr[15:10] == 5'd18);
assign csrbank17_re = interface17_bank_bus_re;
assign csrbank17_ev_soft0_r = interface17_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank17_ev_soft0_re <= 1'd0;
    csrbank17_ev_soft0_we <= 1'd0;
    if ((csrbank17_sel & (interface17_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank17_ev_soft0_re <= interface17_bank_bus_we;
        csrbank17_ev_soft0_we <= csrbank17_re;
    end
end
assign csrbank17_ev_edge_triggered0_r = interface17_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank17_ev_edge_triggered0_we <= 1'd0;
    csrbank17_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank17_sel & (interface17_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank17_ev_edge_triggered0_re <= interface17_bank_bus_we;
        csrbank17_ev_edge_triggered0_we <= csrbank17_re;
    end
end
assign csrbank17_ev_polarity0_r = interface17_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank17_ev_polarity0_we <= 1'd0;
    csrbank17_ev_polarity0_re <= 1'd0;
    if ((csrbank17_sel & (interface17_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank17_ev_polarity0_re <= interface17_bank_bus_we;
        csrbank17_ev_polarity0_we <= csrbank17_re;
    end
end
assign csrbank17_ev_status_r = interface17_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank17_ev_status_re <= 1'd0;
    csrbank17_ev_status_we <= 1'd0;
    if ((csrbank17_sel & (interface17_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank17_ev_status_re <= interface17_bank_bus_we;
        csrbank17_ev_status_we <= csrbank17_re;
    end
end
assign csrbank17_ev_pending_r = interface17_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank17_ev_pending_we <= 1'd0;
    csrbank17_ev_pending_re <= 1'd0;
    if ((csrbank17_sel & (interface17_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank17_ev_pending_re <= interface17_bank_bus_we;
        csrbank17_ev_pending_we <= csrbank17_re;
    end
end
assign csrbank17_ev_enable0_r = interface17_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank17_ev_enable0_we <= 1'd0;
    csrbank17_ev_enable0_re <= 1'd0;
    if ((csrbank17_sel & (interface17_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank17_ev_enable0_re <= interface17_bank_bus_we;
        csrbank17_ev_enable0_we <= csrbank17_re;
    end
end
always @(*) begin
    irqarray4_trigger <= 16'd0;
    if (irqarray4_soft_re) begin
        irqarray4_trigger <= irqarray4_soft_storage[15:0];
    end
end
assign csrbank17_ev_soft0_w = irqarray4_soft_storage[15:0];
assign irqarray4_use_edge = irqarray4_edge_triggered_storage[15:0];
assign csrbank17_ev_edge_triggered0_w = irqarray4_edge_triggered_storage[15:0];
assign irqarray4_rising = irqarray4_polarity_storage[15:0];
assign csrbank17_ev_polarity0_w = irqarray4_polarity_storage[15:0];
always @(*) begin
    irqarray4_status_status <= 16'd0;
    irqarray4_status_status[0] <= irqarray4_trng_done_dupe0;
    irqarray4_status_status[1] <= irqarray4_aes_done_dupe0;
    irqarray4_status_status[2] <= irqarray4_pke_done_dupe0;
    irqarray4_status_status[3] <= irqarray4_hash_done_dupe0;
    irqarray4_status_status[4] <= irqarray4_alu_done_dupe0;
    irqarray4_status_status[5] <= irqarray4_sdma_ichdone_dupe0;
    irqarray4_status_status[6] <= irqarray4_sdma_schdone_dupe0;
    irqarray4_status_status[7] <= irqarray4_sdma_xchdone_dupe0;
    irqarray4_status_status[8] <= irqarray4_nc_b4s80;
    irqarray4_status_status[9] <= irqarray4_nc_b4s90;
    irqarray4_status_status[10] <= irqarray4_nc_b4s100;
    irqarray4_status_status[11] <= irqarray4_nc_b4s110;
    irqarray4_status_status[12] <= irqarray4_nc_b4s120;
    irqarray4_status_status[13] <= irqarray4_nc_b4s130;
    irqarray4_status_status[14] <= irqarray4_nc_b4s140;
    irqarray4_status_status[15] <= irqarray4_nc_b4s150;
end
assign csrbank17_ev_status_w = irqarray4_status_status[15:0];
assign irqarray4_status_we = csrbank17_ev_status_we;
always @(*) begin
    irqarray4_pending_status <= 16'd0;
    irqarray4_pending_status[0] <= irqarray4_trng_done_dupe1;
    irqarray4_pending_status[1] <= irqarray4_aes_done_dupe1;
    irqarray4_pending_status[2] <= irqarray4_pke_done_dupe1;
    irqarray4_pending_status[3] <= irqarray4_hash_done_dupe1;
    irqarray4_pending_status[4] <= irqarray4_alu_done_dupe1;
    irqarray4_pending_status[5] <= irqarray4_sdma_ichdone_dupe1;
    irqarray4_pending_status[6] <= irqarray4_sdma_schdone_dupe1;
    irqarray4_pending_status[7] <= irqarray4_sdma_xchdone_dupe1;
    irqarray4_pending_status[8] <= irqarray4_nc_b4s81;
    irqarray4_pending_status[9] <= irqarray4_nc_b4s91;
    irqarray4_pending_status[10] <= irqarray4_nc_b4s101;
    irqarray4_pending_status[11] <= irqarray4_nc_b4s111;
    irqarray4_pending_status[12] <= irqarray4_nc_b4s121;
    irqarray4_pending_status[13] <= irqarray4_nc_b4s131;
    irqarray4_pending_status[14] <= irqarray4_nc_b4s141;
    irqarray4_pending_status[15] <= irqarray4_nc_b4s151;
end
assign csrbank17_ev_pending_w = irqarray4_pending_status[15:0];
assign irqarray4_pending_we = csrbank17_ev_pending_we;
assign irqarray4_trng_done_dupe2 = irqarray4_enable_storage[0];
assign irqarray4_aes_done_dupe2 = irqarray4_enable_storage[1];
assign irqarray4_pke_done_dupe2 = irqarray4_enable_storage[2];
assign irqarray4_hash_done_dupe2 = irqarray4_enable_storage[3];
assign irqarray4_alu_done_dupe2 = irqarray4_enable_storage[4];
assign irqarray4_sdma_ichdone_dupe2 = irqarray4_enable_storage[5];
assign irqarray4_sdma_schdone_dupe2 = irqarray4_enable_storage[6];
assign irqarray4_sdma_xchdone_dupe2 = irqarray4_enable_storage[7];
assign irqarray4_nc_b4s82 = irqarray4_enable_storage[8];
assign irqarray4_nc_b4s92 = irqarray4_enable_storage[9];
assign irqarray4_nc_b4s102 = irqarray4_enable_storage[10];
assign irqarray4_nc_b4s112 = irqarray4_enable_storage[11];
assign irqarray4_nc_b4s122 = irqarray4_enable_storage[12];
assign irqarray4_nc_b4s132 = irqarray4_enable_storage[13];
assign irqarray4_nc_b4s142 = irqarray4_enable_storage[14];
assign irqarray4_nc_b4s152 = irqarray4_enable_storage[15];
assign csrbank17_ev_enable0_w = irqarray4_enable_storage[15:0];
assign csrbank18_sel = (interface18_bank_bus_adr[15:10] == 5'd19);
assign csrbank18_re = interface18_bank_bus_re;
assign csrbank18_ev_soft0_r = interface18_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank18_ev_soft0_re <= 1'd0;
    csrbank18_ev_soft0_we <= 1'd0;
    if ((csrbank18_sel & (interface18_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank18_ev_soft0_re <= interface18_bank_bus_we;
        csrbank18_ev_soft0_we <= csrbank18_re;
    end
end
assign csrbank18_ev_edge_triggered0_r = interface18_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank18_ev_edge_triggered0_we <= 1'd0;
    csrbank18_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank18_sel & (interface18_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank18_ev_edge_triggered0_re <= interface18_bank_bus_we;
        csrbank18_ev_edge_triggered0_we <= csrbank18_re;
    end
end
assign csrbank18_ev_polarity0_r = interface18_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank18_ev_polarity0_we <= 1'd0;
    csrbank18_ev_polarity0_re <= 1'd0;
    if ((csrbank18_sel & (interface18_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank18_ev_polarity0_re <= interface18_bank_bus_we;
        csrbank18_ev_polarity0_we <= csrbank18_re;
    end
end
assign csrbank18_ev_status_r = interface18_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank18_ev_status_re <= 1'd0;
    csrbank18_ev_status_we <= 1'd0;
    if ((csrbank18_sel & (interface18_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank18_ev_status_re <= interface18_bank_bus_we;
        csrbank18_ev_status_we <= csrbank18_re;
    end
end
assign csrbank18_ev_pending_r = interface18_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank18_ev_pending_we <= 1'd0;
    csrbank18_ev_pending_re <= 1'd0;
    if ((csrbank18_sel & (interface18_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank18_ev_pending_re <= interface18_bank_bus_we;
        csrbank18_ev_pending_we <= csrbank18_re;
    end
end
assign csrbank18_ev_enable0_r = interface18_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank18_ev_enable0_we <= 1'd0;
    csrbank18_ev_enable0_re <= 1'd0;
    if ((csrbank18_sel & (interface18_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank18_ev_enable0_re <= interface18_bank_bus_we;
        csrbank18_ev_enable0_we <= csrbank18_re;
    end
end
always @(*) begin
    irqarray5_trigger <= 16'd0;
    if (irqarray5_soft_re) begin
        irqarray5_trigger <= irqarray5_soft_storage[15:0];
    end
end
assign csrbank18_ev_soft0_w = irqarray5_soft_storage[15:0];
assign irqarray5_use_edge = irqarray5_edge_triggered_storage[15:0];
assign csrbank18_ev_edge_triggered0_w = irqarray5_edge_triggered_storage[15:0];
assign irqarray5_rising = irqarray5_polarity_storage[15:0];
assign csrbank18_ev_polarity0_w = irqarray5_polarity_storage[15:0];
always @(*) begin
    irqarray5_status_status <= 16'd0;
    irqarray5_status_status[0] <= irqarray5_uart0_rx0;
    irqarray5_status_status[1] <= irqarray5_uart0_tx0;
    irqarray5_status_status[2] <= irqarray5_uart0_rx_char0;
    irqarray5_status_status[3] <= irqarray5_uart0_err0;
    irqarray5_status_status[4] <= irqarray5_uart1_rx0;
    irqarray5_status_status[5] <= irqarray5_uart1_tx0;
    irqarray5_status_status[6] <= irqarray5_uart1_rx_char0;
    irqarray5_status_status[7] <= irqarray5_uart1_err0;
    irqarray5_status_status[8] <= irqarray5_uart2_rx0;
    irqarray5_status_status[9] <= irqarray5_uart2_tx0;
    irqarray5_status_status[10] <= irqarray5_uart2_rx_char0;
    irqarray5_status_status[11] <= irqarray5_uart2_err0;
    irqarray5_status_status[12] <= irqarray5_uart3_rx0;
    irqarray5_status_status[13] <= irqarray5_uart3_tx0;
    irqarray5_status_status[14] <= irqarray5_uart3_rx_char0;
    irqarray5_status_status[15] <= irqarray5_uart3_err0;
end
assign csrbank18_ev_status_w = irqarray5_status_status[15:0];
assign irqarray5_status_we = csrbank18_ev_status_we;
always @(*) begin
    irqarray5_pending_status <= 16'd0;
    irqarray5_pending_status[0] <= irqarray5_uart0_rx1;
    irqarray5_pending_status[1] <= irqarray5_uart0_tx1;
    irqarray5_pending_status[2] <= irqarray5_uart0_rx_char1;
    irqarray5_pending_status[3] <= irqarray5_uart0_err1;
    irqarray5_pending_status[4] <= irqarray5_uart1_rx1;
    irqarray5_pending_status[5] <= irqarray5_uart1_tx1;
    irqarray5_pending_status[6] <= irqarray5_uart1_rx_char1;
    irqarray5_pending_status[7] <= irqarray5_uart1_err1;
    irqarray5_pending_status[8] <= irqarray5_uart2_rx1;
    irqarray5_pending_status[9] <= irqarray5_uart2_tx1;
    irqarray5_pending_status[10] <= irqarray5_uart2_rx_char1;
    irqarray5_pending_status[11] <= irqarray5_uart2_err1;
    irqarray5_pending_status[12] <= irqarray5_uart3_rx1;
    irqarray5_pending_status[13] <= irqarray5_uart3_tx1;
    irqarray5_pending_status[14] <= irqarray5_uart3_rx_char1;
    irqarray5_pending_status[15] <= irqarray5_uart3_err1;
end
assign csrbank18_ev_pending_w = irqarray5_pending_status[15:0];
assign irqarray5_pending_we = csrbank18_ev_pending_we;
assign irqarray5_uart0_rx2 = irqarray5_enable_storage[0];
assign irqarray5_uart0_tx2 = irqarray5_enable_storage[1];
assign irqarray5_uart0_rx_char2 = irqarray5_enable_storage[2];
assign irqarray5_uart0_err2 = irqarray5_enable_storage[3];
assign irqarray5_uart1_rx2 = irqarray5_enable_storage[4];
assign irqarray5_uart1_tx2 = irqarray5_enable_storage[5];
assign irqarray5_uart1_rx_char2 = irqarray5_enable_storage[6];
assign irqarray5_uart1_err2 = irqarray5_enable_storage[7];
assign irqarray5_uart2_rx2 = irqarray5_enable_storage[8];
assign irqarray5_uart2_tx2 = irqarray5_enable_storage[9];
assign irqarray5_uart2_rx_char2 = irqarray5_enable_storage[10];
assign irqarray5_uart2_err2 = irqarray5_enable_storage[11];
assign irqarray5_uart3_rx2 = irqarray5_enable_storage[12];
assign irqarray5_uart3_tx2 = irqarray5_enable_storage[13];
assign irqarray5_uart3_rx_char2 = irqarray5_enable_storage[14];
assign irqarray5_uart3_err2 = irqarray5_enable_storage[15];
assign csrbank18_ev_enable0_w = irqarray5_enable_storage[15:0];
assign csrbank19_sel = (interface19_bank_bus_adr[15:10] == 5'd20);
assign csrbank19_re = interface19_bank_bus_re;
assign csrbank19_ev_soft0_r = interface19_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank19_ev_soft0_re <= 1'd0;
    csrbank19_ev_soft0_we <= 1'd0;
    if ((csrbank19_sel & (interface19_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank19_ev_soft0_re <= interface19_bank_bus_we;
        csrbank19_ev_soft0_we <= csrbank19_re;
    end
end
assign csrbank19_ev_edge_triggered0_r = interface19_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank19_ev_edge_triggered0_we <= 1'd0;
    csrbank19_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank19_sel & (interface19_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank19_ev_edge_triggered0_re <= interface19_bank_bus_we;
        csrbank19_ev_edge_triggered0_we <= csrbank19_re;
    end
end
assign csrbank19_ev_polarity0_r = interface19_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank19_ev_polarity0_we <= 1'd0;
    csrbank19_ev_polarity0_re <= 1'd0;
    if ((csrbank19_sel & (interface19_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank19_ev_polarity0_re <= interface19_bank_bus_we;
        csrbank19_ev_polarity0_we <= csrbank19_re;
    end
end
assign csrbank19_ev_status_r = interface19_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank19_ev_status_re <= 1'd0;
    csrbank19_ev_status_we <= 1'd0;
    if ((csrbank19_sel & (interface19_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank19_ev_status_re <= interface19_bank_bus_we;
        csrbank19_ev_status_we <= csrbank19_re;
    end
end
assign csrbank19_ev_pending_r = interface19_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank19_ev_pending_we <= 1'd0;
    csrbank19_ev_pending_re <= 1'd0;
    if ((csrbank19_sel & (interface19_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank19_ev_pending_re <= interface19_bank_bus_we;
        csrbank19_ev_pending_we <= csrbank19_re;
    end
end
assign csrbank19_ev_enable0_r = interface19_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank19_ev_enable0_we <= 1'd0;
    csrbank19_ev_enable0_re <= 1'd0;
    if ((csrbank19_sel & (interface19_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank19_ev_enable0_re <= interface19_bank_bus_we;
        csrbank19_ev_enable0_we <= csrbank19_re;
    end
end
always @(*) begin
    irqarray6_trigger <= 16'd0;
    if (irqarray6_soft_re) begin
        irqarray6_trigger <= irqarray6_soft_storage[15:0];
    end
end
assign csrbank19_ev_soft0_w = irqarray6_soft_storage[15:0];
assign irqarray6_use_edge = irqarray6_edge_triggered_storage[15:0];
assign csrbank19_ev_edge_triggered0_w = irqarray6_edge_triggered_storage[15:0];
assign irqarray6_rising = irqarray6_polarity_storage[15:0];
assign csrbank19_ev_polarity0_w = irqarray6_polarity_storage[15:0];
always @(*) begin
    irqarray6_status_status <= 16'd0;
    irqarray6_status_status[0] <= irqarray6_spim0_rx0;
    irqarray6_status_status[1] <= irqarray6_spim0_tx0;
    irqarray6_status_status[2] <= irqarray6_spim0_cmd0;
    irqarray6_status_status[3] <= irqarray6_spim0_eot0;
    irqarray6_status_status[4] <= irqarray6_spim1_rx0;
    irqarray6_status_status[5] <= irqarray6_spim1_tx0;
    irqarray6_status_status[6] <= irqarray6_spim1_cmd0;
    irqarray6_status_status[7] <= irqarray6_spim1_eot0;
    irqarray6_status_status[8] <= irqarray6_spim2_rx0;
    irqarray6_status_status[9] <= irqarray6_spim2_tx0;
    irqarray6_status_status[10] <= irqarray6_spim2_cmd0;
    irqarray6_status_status[11] <= irqarray6_spim2_eot0;
    irqarray6_status_status[12] <= irqarray6_spim3_rx0;
    irqarray6_status_status[13] <= irqarray6_spim3_tx0;
    irqarray6_status_status[14] <= irqarray6_spim3_cmd0;
    irqarray6_status_status[15] <= irqarray6_spim3_eot0;
end
assign csrbank19_ev_status_w = irqarray6_status_status[15:0];
assign irqarray6_status_we = csrbank19_ev_status_we;
always @(*) begin
    irqarray6_pending_status <= 16'd0;
    irqarray6_pending_status[0] <= irqarray6_spim0_rx1;
    irqarray6_pending_status[1] <= irqarray6_spim0_tx1;
    irqarray6_pending_status[2] <= irqarray6_spim0_cmd1;
    irqarray6_pending_status[3] <= irqarray6_spim0_eot1;
    irqarray6_pending_status[4] <= irqarray6_spim1_rx1;
    irqarray6_pending_status[5] <= irqarray6_spim1_tx1;
    irqarray6_pending_status[6] <= irqarray6_spim1_cmd1;
    irqarray6_pending_status[7] <= irqarray6_spim1_eot1;
    irqarray6_pending_status[8] <= irqarray6_spim2_rx1;
    irqarray6_pending_status[9] <= irqarray6_spim2_tx1;
    irqarray6_pending_status[10] <= irqarray6_spim2_cmd1;
    irqarray6_pending_status[11] <= irqarray6_spim2_eot1;
    irqarray6_pending_status[12] <= irqarray6_spim3_rx1;
    irqarray6_pending_status[13] <= irqarray6_spim3_tx1;
    irqarray6_pending_status[14] <= irqarray6_spim3_cmd1;
    irqarray6_pending_status[15] <= irqarray6_spim3_eot1;
end
assign csrbank19_ev_pending_w = irqarray6_pending_status[15:0];
assign irqarray6_pending_we = csrbank19_ev_pending_we;
assign irqarray6_spim0_rx2 = irqarray6_enable_storage[0];
assign irqarray6_spim0_tx2 = irqarray6_enable_storage[1];
assign irqarray6_spim0_cmd2 = irqarray6_enable_storage[2];
assign irqarray6_spim0_eot2 = irqarray6_enable_storage[3];
assign irqarray6_spim1_rx2 = irqarray6_enable_storage[4];
assign irqarray6_spim1_tx2 = irqarray6_enable_storage[5];
assign irqarray6_spim1_cmd2 = irqarray6_enable_storage[6];
assign irqarray6_spim1_eot2 = irqarray6_enable_storage[7];
assign irqarray6_spim2_rx2 = irqarray6_enable_storage[8];
assign irqarray6_spim2_tx2 = irqarray6_enable_storage[9];
assign irqarray6_spim2_cmd2 = irqarray6_enable_storage[10];
assign irqarray6_spim2_eot2 = irqarray6_enable_storage[11];
assign irqarray6_spim3_rx2 = irqarray6_enable_storage[12];
assign irqarray6_spim3_tx2 = irqarray6_enable_storage[13];
assign irqarray6_spim3_cmd2 = irqarray6_enable_storage[14];
assign irqarray6_spim3_eot2 = irqarray6_enable_storage[15];
assign csrbank19_ev_enable0_w = irqarray6_enable_storage[15:0];
assign csrbank20_sel = (interface20_bank_bus_adr[15:10] == 5'd21);
assign csrbank20_re = interface20_bank_bus_re;
assign csrbank20_ev_soft0_r = interface20_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank20_ev_soft0_re <= 1'd0;
    csrbank20_ev_soft0_we <= 1'd0;
    if ((csrbank20_sel & (interface20_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank20_ev_soft0_re <= interface20_bank_bus_we;
        csrbank20_ev_soft0_we <= csrbank20_re;
    end
end
assign csrbank20_ev_edge_triggered0_r = interface20_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank20_ev_edge_triggered0_we <= 1'd0;
    csrbank20_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank20_sel & (interface20_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank20_ev_edge_triggered0_re <= interface20_bank_bus_we;
        csrbank20_ev_edge_triggered0_we <= csrbank20_re;
    end
end
assign csrbank20_ev_polarity0_r = interface20_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank20_ev_polarity0_we <= 1'd0;
    csrbank20_ev_polarity0_re <= 1'd0;
    if ((csrbank20_sel & (interface20_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank20_ev_polarity0_re <= interface20_bank_bus_we;
        csrbank20_ev_polarity0_we <= csrbank20_re;
    end
end
assign csrbank20_ev_status_r = interface20_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank20_ev_status_re <= 1'd0;
    csrbank20_ev_status_we <= 1'd0;
    if ((csrbank20_sel & (interface20_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank20_ev_status_re <= interface20_bank_bus_we;
        csrbank20_ev_status_we <= csrbank20_re;
    end
end
assign csrbank20_ev_pending_r = interface20_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank20_ev_pending_we <= 1'd0;
    csrbank20_ev_pending_re <= 1'd0;
    if ((csrbank20_sel & (interface20_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank20_ev_pending_re <= interface20_bank_bus_we;
        csrbank20_ev_pending_we <= csrbank20_re;
    end
end
assign csrbank20_ev_enable0_r = interface20_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank20_ev_enable0_we <= 1'd0;
    csrbank20_ev_enable0_re <= 1'd0;
    if ((csrbank20_sel & (interface20_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank20_ev_enable0_re <= interface20_bank_bus_we;
        csrbank20_ev_enable0_we <= csrbank20_re;
    end
end
always @(*) begin
    irqarray7_trigger <= 16'd0;
    if (irqarray7_soft_re) begin
        irqarray7_trigger <= irqarray7_soft_storage[15:0];
    end
end
assign csrbank20_ev_soft0_w = irqarray7_soft_storage[15:0];
assign irqarray7_use_edge = irqarray7_edge_triggered_storage[15:0];
assign csrbank20_ev_edge_triggered0_w = irqarray7_edge_triggered_storage[15:0];
assign irqarray7_rising = irqarray7_polarity_storage[15:0];
assign csrbank20_ev_polarity0_w = irqarray7_polarity_storage[15:0];
always @(*) begin
    irqarray7_status_status <= 16'd0;
    irqarray7_status_status[0] <= irqarray7_i2c0_rx0;
    irqarray7_status_status[1] <= irqarray7_i2c0_tx0;
    irqarray7_status_status[2] <= irqarray7_i2c0_cmd0;
    irqarray7_status_status[3] <= irqarray7_i2c0_eot0;
    irqarray7_status_status[4] <= irqarray7_i2c1_rx0;
    irqarray7_status_status[5] <= irqarray7_i2c1_tx0;
    irqarray7_status_status[6] <= irqarray7_i2c1_cmd0;
    irqarray7_status_status[7] <= irqarray7_i2c1_eot0;
    irqarray7_status_status[8] <= irqarray7_i2c2_rx0;
    irqarray7_status_status[9] <= irqarray7_i2c2_tx0;
    irqarray7_status_status[10] <= irqarray7_i2c2_cmd0;
    irqarray7_status_status[11] <= irqarray7_i2c2_eot0;
    irqarray7_status_status[12] <= irqarray7_i2c3_rx0;
    irqarray7_status_status[13] <= irqarray7_i2c3_tx0;
    irqarray7_status_status[14] <= irqarray7_i2c3_cmd0;
    irqarray7_status_status[15] <= irqarray7_i2c3_eot0;
end
assign csrbank20_ev_status_w = irqarray7_status_status[15:0];
assign irqarray7_status_we = csrbank20_ev_status_we;
always @(*) begin
    irqarray7_pending_status <= 16'd0;
    irqarray7_pending_status[0] <= irqarray7_i2c0_rx1;
    irqarray7_pending_status[1] <= irqarray7_i2c0_tx1;
    irqarray7_pending_status[2] <= irqarray7_i2c0_cmd1;
    irqarray7_pending_status[3] <= irqarray7_i2c0_eot1;
    irqarray7_pending_status[4] <= irqarray7_i2c1_rx1;
    irqarray7_pending_status[5] <= irqarray7_i2c1_tx1;
    irqarray7_pending_status[6] <= irqarray7_i2c1_cmd1;
    irqarray7_pending_status[7] <= irqarray7_i2c1_eot1;
    irqarray7_pending_status[8] <= irqarray7_i2c2_rx1;
    irqarray7_pending_status[9] <= irqarray7_i2c2_tx1;
    irqarray7_pending_status[10] <= irqarray7_i2c2_cmd1;
    irqarray7_pending_status[11] <= irqarray7_i2c2_eot1;
    irqarray7_pending_status[12] <= irqarray7_i2c3_rx1;
    irqarray7_pending_status[13] <= irqarray7_i2c3_tx1;
    irqarray7_pending_status[14] <= irqarray7_i2c3_cmd1;
    irqarray7_pending_status[15] <= irqarray7_i2c3_eot1;
end
assign csrbank20_ev_pending_w = irqarray7_pending_status[15:0];
assign irqarray7_pending_we = csrbank20_ev_pending_we;
assign irqarray7_i2c0_rx2 = irqarray7_enable_storage[0];
assign irqarray7_i2c0_tx2 = irqarray7_enable_storage[1];
assign irqarray7_i2c0_cmd2 = irqarray7_enable_storage[2];
assign irqarray7_i2c0_eot2 = irqarray7_enable_storage[3];
assign irqarray7_i2c1_rx2 = irqarray7_enable_storage[4];
assign irqarray7_i2c1_tx2 = irqarray7_enable_storage[5];
assign irqarray7_i2c1_cmd2 = irqarray7_enable_storage[6];
assign irqarray7_i2c1_eot2 = irqarray7_enable_storage[7];
assign irqarray7_i2c2_rx2 = irqarray7_enable_storage[8];
assign irqarray7_i2c2_tx2 = irqarray7_enable_storage[9];
assign irqarray7_i2c2_cmd2 = irqarray7_enable_storage[10];
assign irqarray7_i2c2_eot2 = irqarray7_enable_storage[11];
assign irqarray7_i2c3_rx2 = irqarray7_enable_storage[12];
assign irqarray7_i2c3_tx2 = irqarray7_enable_storage[13];
assign irqarray7_i2c3_cmd2 = irqarray7_enable_storage[14];
assign irqarray7_i2c3_eot2 = irqarray7_enable_storage[15];
assign csrbank20_ev_enable0_w = irqarray7_enable_storage[15:0];
assign csrbank21_sel = (interface21_bank_bus_adr[15:10] == 5'd22);
assign csrbank21_re = interface21_bank_bus_re;
assign csrbank21_ev_soft0_r = interface21_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank21_ev_soft0_re <= 1'd0;
    csrbank21_ev_soft0_we <= 1'd0;
    if ((csrbank21_sel & (interface21_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank21_ev_soft0_re <= interface21_bank_bus_we;
        csrbank21_ev_soft0_we <= csrbank21_re;
    end
end
assign csrbank21_ev_edge_triggered0_r = interface21_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank21_ev_edge_triggered0_we <= 1'd0;
    csrbank21_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank21_sel & (interface21_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank21_ev_edge_triggered0_re <= interface21_bank_bus_we;
        csrbank21_ev_edge_triggered0_we <= csrbank21_re;
    end
end
assign csrbank21_ev_polarity0_r = interface21_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank21_ev_polarity0_we <= 1'd0;
    csrbank21_ev_polarity0_re <= 1'd0;
    if ((csrbank21_sel & (interface21_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank21_ev_polarity0_re <= interface21_bank_bus_we;
        csrbank21_ev_polarity0_we <= csrbank21_re;
    end
end
assign csrbank21_ev_status_r = interface21_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank21_ev_status_re <= 1'd0;
    csrbank21_ev_status_we <= 1'd0;
    if ((csrbank21_sel & (interface21_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank21_ev_status_re <= interface21_bank_bus_we;
        csrbank21_ev_status_we <= csrbank21_re;
    end
end
assign csrbank21_ev_pending_r = interface21_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank21_ev_pending_we <= 1'd0;
    csrbank21_ev_pending_re <= 1'd0;
    if ((csrbank21_sel & (interface21_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank21_ev_pending_re <= interface21_bank_bus_we;
        csrbank21_ev_pending_we <= csrbank21_re;
    end
end
assign csrbank21_ev_enable0_r = interface21_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank21_ev_enable0_we <= 1'd0;
    csrbank21_ev_enable0_re <= 1'd0;
    if ((csrbank21_sel & (interface21_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank21_ev_enable0_re <= interface21_bank_bus_we;
        csrbank21_ev_enable0_we <= csrbank21_re;
    end
end
always @(*) begin
    irqarray8_trigger <= 16'd0;
    if (irqarray8_soft_re) begin
        irqarray8_trigger <= irqarray8_soft_storage[15:0];
    end
end
assign csrbank21_ev_soft0_w = irqarray8_soft_storage[15:0];
assign irqarray8_use_edge = irqarray8_edge_triggered_storage[15:0];
assign csrbank21_ev_edge_triggered0_w = irqarray8_edge_triggered_storage[15:0];
assign irqarray8_rising = irqarray8_polarity_storage[15:0];
assign csrbank21_ev_polarity0_w = irqarray8_polarity_storage[15:0];
always @(*) begin
    irqarray8_status_status <= 16'd0;
    irqarray8_status_status[0] <= irqarray8_sdio_rx0;
    irqarray8_status_status[1] <= irqarray8_sdio_tx0;
    irqarray8_status_status[2] <= irqarray8_sdio_eot0;
    irqarray8_status_status[3] <= irqarray8_sdio_err0;
    irqarray8_status_status[4] <= irqarray8_i2s_rx0;
    irqarray8_status_status[5] <= irqarray8_i2s_tx0;
    irqarray8_status_status[6] <= irqarray8_nc_b8s60;
    irqarray8_status_status[7] <= irqarray8_nc_b8s70;
    irqarray8_status_status[8] <= irqarray8_cam_rx0;
    irqarray8_status_status[9] <= irqarray8_adc_rx0;
    irqarray8_status_status[10] <= irqarray8_nc_b8s100;
    irqarray8_status_status[11] <= irqarray8_nc_b8s110;
    irqarray8_status_status[12] <= irqarray8_filter_eot0;
    irqarray8_status_status[13] <= irqarray8_filter_act0;
    irqarray8_status_status[14] <= irqarray8_nc_b8s140;
    irqarray8_status_status[15] <= irqarray8_nc_b8s150;
end
assign csrbank21_ev_status_w = irqarray8_status_status[15:0];
assign irqarray8_status_we = csrbank21_ev_status_we;
always @(*) begin
    irqarray8_pending_status <= 16'd0;
    irqarray8_pending_status[0] <= irqarray8_sdio_rx1;
    irqarray8_pending_status[1] <= irqarray8_sdio_tx1;
    irqarray8_pending_status[2] <= irqarray8_sdio_eot1;
    irqarray8_pending_status[3] <= irqarray8_sdio_err1;
    irqarray8_pending_status[4] <= irqarray8_i2s_rx1;
    irqarray8_pending_status[5] <= irqarray8_i2s_tx1;
    irqarray8_pending_status[6] <= irqarray8_nc_b8s61;
    irqarray8_pending_status[7] <= irqarray8_nc_b8s71;
    irqarray8_pending_status[8] <= irqarray8_cam_rx1;
    irqarray8_pending_status[9] <= irqarray8_adc_rx1;
    irqarray8_pending_status[10] <= irqarray8_nc_b8s101;
    irqarray8_pending_status[11] <= irqarray8_nc_b8s111;
    irqarray8_pending_status[12] <= irqarray8_filter_eot1;
    irqarray8_pending_status[13] <= irqarray8_filter_act1;
    irqarray8_pending_status[14] <= irqarray8_nc_b8s141;
    irqarray8_pending_status[15] <= irqarray8_nc_b8s151;
end
assign csrbank21_ev_pending_w = irqarray8_pending_status[15:0];
assign irqarray8_pending_we = csrbank21_ev_pending_we;
assign irqarray8_sdio_rx2 = irqarray8_enable_storage[0];
assign irqarray8_sdio_tx2 = irqarray8_enable_storage[1];
assign irqarray8_sdio_eot2 = irqarray8_enable_storage[2];
assign irqarray8_sdio_err2 = irqarray8_enable_storage[3];
assign irqarray8_i2s_rx2 = irqarray8_enable_storage[4];
assign irqarray8_i2s_tx2 = irqarray8_enable_storage[5];
assign irqarray8_nc_b8s62 = irqarray8_enable_storage[6];
assign irqarray8_nc_b8s72 = irqarray8_enable_storage[7];
assign irqarray8_cam_rx2 = irqarray8_enable_storage[8];
assign irqarray8_adc_rx2 = irqarray8_enable_storage[9];
assign irqarray8_nc_b8s102 = irqarray8_enable_storage[10];
assign irqarray8_nc_b8s112 = irqarray8_enable_storage[11];
assign irqarray8_filter_eot2 = irqarray8_enable_storage[12];
assign irqarray8_filter_act2 = irqarray8_enable_storage[13];
assign irqarray8_nc_b8s142 = irqarray8_enable_storage[14];
assign irqarray8_nc_b8s152 = irqarray8_enable_storage[15];
assign csrbank21_ev_enable0_w = irqarray8_enable_storage[15:0];
assign csrbank22_sel = (interface22_bank_bus_adr[15:10] == 5'd23);
assign csrbank22_re = interface22_bank_bus_re;
assign csrbank22_ev_soft0_r = interface22_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank22_ev_soft0_re <= 1'd0;
    csrbank22_ev_soft0_we <= 1'd0;
    if ((csrbank22_sel & (interface22_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank22_ev_soft0_re <= interface22_bank_bus_we;
        csrbank22_ev_soft0_we <= csrbank22_re;
    end
end
assign csrbank22_ev_edge_triggered0_r = interface22_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank22_ev_edge_triggered0_we <= 1'd0;
    csrbank22_ev_edge_triggered0_re <= 1'd0;
    if ((csrbank22_sel & (interface22_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank22_ev_edge_triggered0_re <= interface22_bank_bus_we;
        csrbank22_ev_edge_triggered0_we <= csrbank22_re;
    end
end
assign csrbank22_ev_polarity0_r = interface22_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank22_ev_polarity0_we <= 1'd0;
    csrbank22_ev_polarity0_re <= 1'd0;
    if ((csrbank22_sel & (interface22_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank22_ev_polarity0_re <= interface22_bank_bus_we;
        csrbank22_ev_polarity0_we <= csrbank22_re;
    end
end
assign csrbank22_ev_status_r = interface22_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank22_ev_status_re <= 1'd0;
    csrbank22_ev_status_we <= 1'd0;
    if ((csrbank22_sel & (interface22_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank22_ev_status_re <= interface22_bank_bus_we;
        csrbank22_ev_status_we <= csrbank22_re;
    end
end
assign csrbank22_ev_pending_r = interface22_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank22_ev_pending_we <= 1'd0;
    csrbank22_ev_pending_re <= 1'd0;
    if ((csrbank22_sel & (interface22_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank22_ev_pending_re <= interface22_bank_bus_we;
        csrbank22_ev_pending_we <= csrbank22_re;
    end
end
assign csrbank22_ev_enable0_r = interface22_bank_bus_dat_w[15:0];
always @(*) begin
    csrbank22_ev_enable0_we <= 1'd0;
    csrbank22_ev_enable0_re <= 1'd0;
    if ((csrbank22_sel & (interface22_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank22_ev_enable0_re <= interface22_bank_bus_we;
        csrbank22_ev_enable0_we <= csrbank22_re;
    end
end
always @(*) begin
    irqarray9_trigger <= 16'd0;
    if (irqarray9_soft_re) begin
        irqarray9_trigger <= irqarray9_soft_storage[15:0];
    end
end
assign csrbank22_ev_soft0_w = irqarray9_soft_storage[15:0];
assign irqarray9_use_edge = irqarray9_edge_triggered_storage[15:0];
assign csrbank22_ev_edge_triggered0_w = irqarray9_edge_triggered_storage[15:0];
assign irqarray9_rising = irqarray9_polarity_storage[15:0];
assign csrbank22_ev_polarity0_w = irqarray9_polarity_storage[15:0];
always @(*) begin
    irqarray9_status_status <= 16'd0;
    irqarray9_status_status[0] <= irqarray9_scif_rx0;
    irqarray9_status_status[1] <= irqarray9_scif_tx0;
    irqarray9_status_status[2] <= irqarray9_scif_rx_char0;
    irqarray9_status_status[3] <= irqarray9_scif_err0;
    irqarray9_status_status[4] <= irqarray9_spis0_rx0;
    irqarray9_status_status[5] <= irqarray9_spis0_tx0;
    irqarray9_status_status[6] <= irqarray9_spis0_eot0;
    irqarray9_status_status[7] <= irqarray9_nc_b9s70;
    irqarray9_status_status[8] <= irqarray9_spis1_rx0;
    irqarray9_status_status[9] <= irqarray9_spis1_tx0;
    irqarray9_status_status[10] <= irqarray9_spis1_eot0;
    irqarray9_status_status[11] <= irqarray9_nc_b9s110;
    irqarray9_status_status[12] <= irqarray9_pwm0_ev0;
    irqarray9_status_status[13] <= irqarray9_pwm1_ev0;
    irqarray9_status_status[14] <= irqarray9_pwm2_ev0;
    irqarray9_status_status[15] <= irqarray9_pwm3_ev0;
end
assign csrbank22_ev_status_w = irqarray9_status_status[15:0];
assign irqarray9_status_we = csrbank22_ev_status_we;
always @(*) begin
    irqarray9_pending_status <= 16'd0;
    irqarray9_pending_status[0] <= irqarray9_scif_rx1;
    irqarray9_pending_status[1] <= irqarray9_scif_tx1;
    irqarray9_pending_status[2] <= irqarray9_scif_rx_char1;
    irqarray9_pending_status[3] <= irqarray9_scif_err1;
    irqarray9_pending_status[4] <= irqarray9_spis0_rx1;
    irqarray9_pending_status[5] <= irqarray9_spis0_tx1;
    irqarray9_pending_status[6] <= irqarray9_spis0_eot1;
    irqarray9_pending_status[7] <= irqarray9_nc_b9s71;
    irqarray9_pending_status[8] <= irqarray9_spis1_rx1;
    irqarray9_pending_status[9] <= irqarray9_spis1_tx1;
    irqarray9_pending_status[10] <= irqarray9_spis1_eot1;
    irqarray9_pending_status[11] <= irqarray9_nc_b9s111;
    irqarray9_pending_status[12] <= irqarray9_pwm0_ev1;
    irqarray9_pending_status[13] <= irqarray9_pwm1_ev1;
    irqarray9_pending_status[14] <= irqarray9_pwm2_ev1;
    irqarray9_pending_status[15] <= irqarray9_pwm3_ev1;
end
assign csrbank22_ev_pending_w = irqarray9_pending_status[15:0];
assign irqarray9_pending_we = csrbank22_ev_pending_we;
assign irqarray9_scif_rx2 = irqarray9_enable_storage[0];
assign irqarray9_scif_tx2 = irqarray9_enable_storage[1];
assign irqarray9_scif_rx_char2 = irqarray9_enable_storage[2];
assign irqarray9_scif_err2 = irqarray9_enable_storage[3];
assign irqarray9_spis0_rx2 = irqarray9_enable_storage[4];
assign irqarray9_spis0_tx2 = irqarray9_enable_storage[5];
assign irqarray9_spis0_eot2 = irqarray9_enable_storage[6];
assign irqarray9_nc_b9s72 = irqarray9_enable_storage[7];
assign irqarray9_spis1_rx2 = irqarray9_enable_storage[8];
assign irqarray9_spis1_tx2 = irqarray9_enable_storage[9];
assign irqarray9_spis1_eot2 = irqarray9_enable_storage[10];
assign irqarray9_nc_b9s112 = irqarray9_enable_storage[11];
assign irqarray9_pwm0_ev2 = irqarray9_enable_storage[12];
assign irqarray9_pwm1_ev2 = irqarray9_enable_storage[13];
assign irqarray9_pwm2_ev2 = irqarray9_enable_storage[14];
assign irqarray9_pwm3_ev2 = irqarray9_enable_storage[15];
assign csrbank22_ev_enable0_w = irqarray9_enable_storage[15:0];
assign csrbank23_sel = (interface23_bank_bus_adr[15:10] == 5'd24);
assign csrbank23_re = interface23_bank_bus_re;
assign csrbank23_wdata0_r = interface23_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank23_wdata0_re <= 1'd0;
    csrbank23_wdata0_we <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank23_wdata0_re <= interface23_bank_bus_we;
        csrbank23_wdata0_we <= csrbank23_re;
    end
end
assign csrbank23_rdata_r = interface23_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank23_rdata_we <= 1'd0;
    csrbank23_rdata_re <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank23_rdata_re <= interface23_bank_bus_we;
        csrbank23_rdata_we <= csrbank23_re;
    end
end
assign csrbank23_ev_status_r = interface23_bank_bus_dat_w[3:0];
always @(*) begin
    csrbank23_ev_status_we <= 1'd0;
    csrbank23_ev_status_re <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank23_ev_status_re <= interface23_bank_bus_we;
        csrbank23_ev_status_we <= csrbank23_re;
    end
end
assign csrbank23_ev_pending_r = interface23_bank_bus_dat_w[3:0];
always @(*) begin
    csrbank23_ev_pending_re <= 1'd0;
    csrbank23_ev_pending_we <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank23_ev_pending_re <= interface23_bank_bus_we;
        csrbank23_ev_pending_we <= csrbank23_re;
    end
end
assign csrbank23_ev_enable0_r = interface23_bank_bus_dat_w[3:0];
always @(*) begin
    csrbank23_ev_enable0_re <= 1'd0;
    csrbank23_ev_enable0_we <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank23_ev_enable0_re <= interface23_bank_bus_we;
        csrbank23_ev_enable0_we <= csrbank23_re;
    end
end
assign csrbank23_status_r = interface23_bank_bus_dat_w[25:0];
always @(*) begin
    csrbank23_status_we <= 1'd0;
    csrbank23_status_re <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank23_status_re <= interface23_bank_bus_we;
        csrbank23_status_we <= csrbank23_re;
    end
end
assign csrbank23_control0_r = interface23_bank_bus_dat_w[0];
always @(*) begin
    csrbank23_control0_re <= 1'd0;
    csrbank23_control0_we <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 3'd6))) begin
        csrbank23_control0_re <= interface23_bank_bus_we;
        csrbank23_control0_we <= csrbank23_re;
    end
end
assign csrbank23_done0_r = interface23_bank_bus_dat_w[0];
always @(*) begin
    csrbank23_done0_re <= 1'd0;
    csrbank23_done0_we <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 3'd7))) begin
        csrbank23_done0_re <= interface23_bank_bus_we;
        csrbank23_done0_we <= csrbank23_re;
    end
end
assign csrbank23_loopback0_r = interface23_bank_bus_dat_w[0];
always @(*) begin
    csrbank23_loopback0_we <= 1'd0;
    csrbank23_loopback0_re <= 1'd0;
    if ((csrbank23_sel & (interface23_bank_bus_adr[9:0] == 4'd8))) begin
        csrbank23_loopback0_re <= interface23_bank_bus_we;
        csrbank23_loopback0_we <= csrbank23_re;
    end
end
assign csrbank23_wdata0_w = mailbox_wdata_storage[31:0];
assign csrbank23_rdata_w = mailbox_rdata_status[31:0];
assign mailbox_rdata_we = csrbank23_rdata_we;
always @(*) begin
    mailbox_status_status0 <= 4'd0;
    mailbox_status_status0[0] <= mailbox_available0;
    mailbox_status_status0[1] <= mailbox_abort_init0;
    mailbox_status_status0[2] <= mailbox_abort_done0;
    mailbox_status_status0[3] <= mailbox_error0;
end
assign csrbank23_ev_status_w = mailbox_status_status0[3:0];
assign mailbox_status_we0 = csrbank23_ev_status_we;
always @(*) begin
    mailbox_pending_status <= 4'd0;
    mailbox_pending_status[0] <= mailbox_available1;
    mailbox_pending_status[1] <= mailbox_abort_init1;
    mailbox_pending_status[2] <= mailbox_abort_done1;
    mailbox_pending_status[3] <= mailbox_error1;
end
assign csrbank23_ev_pending_w = mailbox_pending_status[3:0];
assign mailbox_pending_we = csrbank23_ev_pending_we;
assign mailbox_available2 = mailbox_enable_storage[0];
assign mailbox_abort_init2 = mailbox_enable_storage[1];
assign mailbox_abort_done2 = mailbox_enable_storage[2];
assign mailbox_error2 = mailbox_enable_storage[3];
assign csrbank23_ev_enable0_w = mailbox_enable_storage[3:0];
always @(*) begin
    mailbox_status_status1 <= 26'd0;
    mailbox_status_status1[10:0] <= mailbox_rx_words;
    mailbox_status_status1[21:11] <= mailbox_tx_words;
    mailbox_status_status1[22] <= mailbox_abort_in_progress0;
    mailbox_status_status1[23] <= mailbox_abort_ack0;
    mailbox_status_status1[24] <= mailbox_tx_err;
    mailbox_status_status1[25] <= mailbox_rx_err;
end
assign csrbank23_status_w = mailbox_status_status1[25:0];
assign mailbox_status_we1 = csrbank23_status_we;
always @(*) begin
    mailbox_abort <= 1'd0;
    if (mailbox_control_re) begin
        mailbox_abort <= mailbox_control_storage;
    end
end
assign csrbank23_control0_w = mailbox_control_storage;
always @(*) begin
    mailbox_done <= 1'd0;
    if (mailbox_done_re) begin
        mailbox_done <= mailbox_done_storage;
    end
end
assign csrbank23_done0_w = mailbox_done_storage;
assign mailbox_loopback = mailbox_loopback_storage;
assign csrbank23_loopback0_w = mailbox_loopback_storage;
assign csrbank24_sel = (interface24_bank_bus_adr[15:10] == 5'd25);
assign csrbank24_re = interface24_bank_bus_re;
assign csrbank24_wdata0_r = interface24_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank24_wdata0_re <= 1'd0;
    csrbank24_wdata0_we <= 1'd0;
    if ((csrbank24_sel & (interface24_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank24_wdata0_re <= interface24_bank_bus_we;
        csrbank24_wdata0_we <= csrbank24_re;
    end
end
assign csrbank24_rdata_r = interface24_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank24_rdata_we <= 1'd0;
    csrbank24_rdata_re <= 1'd0;
    if ((csrbank24_sel & (interface24_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank24_rdata_re <= interface24_bank_bus_we;
        csrbank24_rdata_we <= csrbank24_re;
    end
end
assign csrbank24_status_r = interface24_bank_bus_dat_w[5:0];
always @(*) begin
    csrbank24_status_we <= 1'd0;
    csrbank24_status_re <= 1'd0;
    if ((csrbank24_sel & (interface24_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank24_status_re <= interface24_bank_bus_we;
        csrbank24_status_we <= csrbank24_re;
    end
end
assign csrbank24_ev_status_r = interface24_bank_bus_dat_w[3:0];
always @(*) begin
    csrbank24_ev_status_re <= 1'd0;
    csrbank24_ev_status_we <= 1'd0;
    if ((csrbank24_sel & (interface24_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank24_ev_status_re <= interface24_bank_bus_we;
        csrbank24_ev_status_we <= csrbank24_re;
    end
end
assign csrbank24_ev_pending_r = interface24_bank_bus_dat_w[3:0];
always @(*) begin
    csrbank24_ev_pending_re <= 1'd0;
    csrbank24_ev_pending_we <= 1'd0;
    if ((csrbank24_sel & (interface24_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank24_ev_pending_re <= interface24_bank_bus_we;
        csrbank24_ev_pending_we <= csrbank24_re;
    end
end
assign csrbank24_ev_enable0_r = interface24_bank_bus_dat_w[3:0];
always @(*) begin
    csrbank24_ev_enable0_we <= 1'd0;
    csrbank24_ev_enable0_re <= 1'd0;
    if ((csrbank24_sel & (interface24_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank24_ev_enable0_re <= interface24_bank_bus_we;
        csrbank24_ev_enable0_we <= csrbank24_re;
    end
end
assign csrbank24_control0_r = interface24_bank_bus_dat_w[0];
always @(*) begin
    csrbank24_control0_re <= 1'd0;
    csrbank24_control0_we <= 1'd0;
    if ((csrbank24_sel & (interface24_bank_bus_adr[9:0] == 3'd6))) begin
        csrbank24_control0_re <= interface24_bank_bus_we;
        csrbank24_control0_we <= csrbank24_re;
    end
end
assign csrbank24_done0_r = interface24_bank_bus_dat_w[0];
always @(*) begin
    csrbank24_done0_we <= 1'd0;
    csrbank24_done0_re <= 1'd0;
    if ((csrbank24_sel & (interface24_bank_bus_adr[9:0] == 3'd7))) begin
        csrbank24_done0_re <= interface24_bank_bus_we;
        csrbank24_done0_we <= csrbank24_re;
    end
end
assign csrbank24_wdata0_w = mb_client_wdata_storage[31:0];
assign csrbank24_rdata_w = mb_client_rdata_status[31:0];
assign mb_client_rdata_we = csrbank24_rdata_we;
always @(*) begin
    mb_client_status_status0 <= 6'd0;
    mb_client_status_status0[0] <= mb_client_rx_avail;
    mb_client_status_status0[1] <= mb_client_tx_free;
    mb_client_status_status0[2] <= mb_client_abort_in_progress0;
    mb_client_status_status0[3] <= mb_client_abort_ack0;
    mb_client_status_status0[4] <= mb_client_tx_err;
    mb_client_status_status0[5] <= mb_client_rx_err;
end
assign csrbank24_status_w = mb_client_status_status0[5:0];
assign mb_client_status_we0 = csrbank24_status_we;
always @(*) begin
    mb_client_status_status1 <= 4'd0;
    mb_client_status_status1[0] <= mb_client_available0;
    mb_client_status_status1[1] <= mb_client_abort_init0;
    mb_client_status_status1[2] <= mb_client_abort_done0;
    mb_client_status_status1[3] <= mb_client_error0;
end
assign csrbank24_ev_status_w = mb_client_status_status1[3:0];
assign mb_client_status_we1 = csrbank24_ev_status_we;
always @(*) begin
    mb_client_pending_status <= 4'd0;
    mb_client_pending_status[0] <= mb_client_available1;
    mb_client_pending_status[1] <= mb_client_abort_init1;
    mb_client_pending_status[2] <= mb_client_abort_done1;
    mb_client_pending_status[3] <= mb_client_error1;
end
assign csrbank24_ev_pending_w = mb_client_pending_status[3:0];
assign mb_client_pending_we = csrbank24_ev_pending_we;
assign mb_client_available2 = mb_client_enable_storage[0];
assign mb_client_abort_init2 = mb_client_enable_storage[1];
assign mb_client_abort_done2 = mb_client_enable_storage[2];
assign mb_client_error2 = mb_client_enable_storage[3];
assign csrbank24_ev_enable0_w = mb_client_enable_storage[3:0];
always @(*) begin
    mb_client_abort <= 1'd0;
    if (mb_client_control_re) begin
        mb_client_abort <= mb_client_control_storage;
    end
end
assign csrbank24_control0_w = mb_client_control_storage;
always @(*) begin
    mb_client_done <= 1'd0;
    if (mb_client_done_re) begin
        mb_client_done <= mb_client_done_storage;
    end
end
assign csrbank24_done0_w = mb_client_done_storage;
assign csrbank25_sel = (interface25_bank_bus_adr[15:10] == 5'd26);
assign csrbank25_re = interface25_bank_bus_re;
assign csrbank25_pc_r = interface25_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank25_pc_re <= 1'd0;
    csrbank25_pc_we <= 1'd0;
    if ((csrbank25_sel & (interface25_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank25_pc_re <= interface25_bank_bus_we;
        csrbank25_pc_we <= csrbank25_re;
    end
end
assign csrbank25_pc_w = status[31:0];
assign we = csrbank25_pc_we;
assign csrbank26_sel = (interface26_bank_bus_adr[15:10] == 1'd1);
assign csrbank26_re = interface26_bank_bus_re;
assign csrbank26_control0_r = interface26_bank_bus_dat_w[1:0];
always @(*) begin
    csrbank26_control0_we <= 1'd0;
    csrbank26_control0_re <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank26_control0_re <= interface26_bank_bus_we;
        csrbank26_control0_we <= csrbank26_re;
    end
end
assign csrbank26_resume_time1_r = interface26_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank26_resume_time1_re <= 1'd0;
    csrbank26_resume_time1_we <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank26_resume_time1_re <= interface26_bank_bus_we;
        csrbank26_resume_time1_we <= csrbank26_re;
    end
end
assign csrbank26_resume_time0_r = interface26_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank26_resume_time0_re <= 1'd0;
    csrbank26_resume_time0_we <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank26_resume_time0_re <= interface26_bank_bus_we;
        csrbank26_resume_time0_we <= csrbank26_re;
    end
end
assign csrbank26_time1_r = interface26_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank26_time1_we <= 1'd0;
    csrbank26_time1_re <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank26_time1_re <= interface26_bank_bus_we;
        csrbank26_time1_we <= csrbank26_re;
    end
end
assign csrbank26_time0_r = interface26_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank26_time0_re <= 1'd0;
    csrbank26_time0_we <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank26_time0_re <= interface26_bank_bus_we;
        csrbank26_time0_we <= csrbank26_re;
    end
end
assign csrbank26_status_r = interface26_bank_bus_dat_w[0];
always @(*) begin
    csrbank26_status_re <= 1'd0;
    csrbank26_status_we <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank26_status_re <= interface26_bank_bus_we;
        csrbank26_status_we <= csrbank26_re;
    end
end
assign csrbank26_state0_r = interface26_bank_bus_dat_w[1:0];
always @(*) begin
    csrbank26_state0_we <= 1'd0;
    csrbank26_state0_re <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 3'd6))) begin
        csrbank26_state0_re <= interface26_bank_bus_we;
        csrbank26_state0_we <= csrbank26_re;
    end
end
assign csrbank26_interrupt0_r = interface26_bank_bus_dat_w[0];
always @(*) begin
    csrbank26_interrupt0_we <= 1'd0;
    csrbank26_interrupt0_re <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 3'd7))) begin
        csrbank26_interrupt0_re <= interface26_bank_bus_we;
        csrbank26_interrupt0_we <= csrbank26_re;
    end
end
assign csrbank26_ev_status_r = interface26_bank_bus_dat_w[0];
always @(*) begin
    csrbank26_ev_status_re <= 1'd0;
    csrbank26_ev_status_we <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 4'd8))) begin
        csrbank26_ev_status_re <= interface26_bank_bus_we;
        csrbank26_ev_status_we <= csrbank26_re;
    end
end
assign csrbank26_ev_pending_r = interface26_bank_bus_dat_w[0];
always @(*) begin
    csrbank26_ev_pending_we <= 1'd0;
    csrbank26_ev_pending_re <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 4'd9))) begin
        csrbank26_ev_pending_re <= interface26_bank_bus_we;
        csrbank26_ev_pending_we <= csrbank26_re;
    end
end
assign csrbank26_ev_enable0_r = interface26_bank_bus_dat_w[0];
always @(*) begin
    csrbank26_ev_enable0_we <= 1'd0;
    csrbank26_ev_enable0_re <= 1'd0;
    if ((csrbank26_sel & (interface26_bank_bus_adr[9:0] == 4'd10))) begin
        csrbank26_ev_enable0_re <= interface26_bank_bus_we;
        csrbank26_ev_enable0_we <= csrbank26_re;
    end
end
assign susres_pause = susres_control_storage[0];
always @(*) begin
    susres_load <= 1'd0;
    if (susres_control_re) begin
        susres_load <= susres_control_storage[1];
    end
end
assign csrbank26_control0_w = susres_control_storage[1:0];
assign csrbank26_resume_time1_w = susres_resume_time_storage[63:32];
assign csrbank26_resume_time0_w = susres_resume_time_storage[31:0];
assign csrbank26_time1_w = susres_time_status[63:32];
assign csrbank26_time0_w = susres_time_status[31:0];
assign susres_time_we = csrbank26_time0_we;
assign susres_status_status0 = susres_paused;
assign csrbank26_status_w = susres_status_status0;
assign susres_status_we0 = csrbank26_status_we;
assign susres_resume0 = susres_state_storage[0];
assign susres_was_forced = susres_state_storage[1];
assign csrbank26_state0_w = susres_state_storage[1:0];
always @(*) begin
    susres_interrupt <= 1'd0;
    if (susres_interrupt_re) begin
        susres_interrupt <= susres_interrupt_storage;
    end
end
assign csrbank26_interrupt0_w = susres_interrupt_storage;
assign susres_status_status1 = susres_soft_int0;
assign csrbank26_ev_status_w = susres_status_status1;
assign susres_status_we1 = csrbank26_ev_status_we;
assign susres_pending_status = susres_soft_int1;
assign csrbank26_ev_pending_w = susres_pending_status;
assign susres_pending_we = csrbank26_ev_pending_we;
assign susres_soft_int2 = susres_enable_storage;
assign csrbank26_ev_enable0_w = susres_enable_storage;
assign csrbank27_sel = (interface27_bank_bus_adr[15:10] == 5'd27);
assign csrbank27_re = interface27_bank_bus_re;
assign csrbank27_control0_r = interface27_bank_bus_dat_w[0];
always @(*) begin
    csrbank27_control0_we <= 1'd0;
    csrbank27_control0_re <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank27_control0_re <= interface27_bank_bus_we;
        csrbank27_control0_we <= csrbank27_re;
    end
end
assign csrbank27_time1_r = interface27_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank27_time1_re <= 1'd0;
    csrbank27_time1_we <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank27_time1_re <= interface27_bank_bus_we;
        csrbank27_time1_we <= csrbank27_re;
    end
end
assign csrbank27_time0_r = interface27_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank27_time0_we <= 1'd0;
    csrbank27_time0_re <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank27_time0_re <= interface27_bank_bus_we;
        csrbank27_time0_we <= csrbank27_re;
    end
end
assign csrbank27_msleep_target1_r = interface27_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank27_msleep_target1_we <= 1'd0;
    csrbank27_msleep_target1_re <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank27_msleep_target1_re <= interface27_bank_bus_we;
        csrbank27_msleep_target1_we <= csrbank27_re;
    end
end
assign csrbank27_msleep_target0_r = interface27_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank27_msleep_target0_re <= 1'd0;
    csrbank27_msleep_target0_we <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank27_msleep_target0_re <= interface27_bank_bus_we;
        csrbank27_msleep_target0_we <= csrbank27_re;
    end
end
assign csrbank27_ev_status_r = interface27_bank_bus_dat_w[0];
always @(*) begin
    csrbank27_ev_status_we <= 1'd0;
    csrbank27_ev_status_re <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank27_ev_status_re <= interface27_bank_bus_we;
        csrbank27_ev_status_we <= csrbank27_re;
    end
end
assign csrbank27_ev_pending_r = interface27_bank_bus_dat_w[0];
always @(*) begin
    csrbank27_ev_pending_we <= 1'd0;
    csrbank27_ev_pending_re <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 3'd6))) begin
        csrbank27_ev_pending_re <= interface27_bank_bus_we;
        csrbank27_ev_pending_we <= csrbank27_re;
    end
end
assign csrbank27_ev_enable0_r = interface27_bank_bus_dat_w[0];
always @(*) begin
    csrbank27_ev_enable0_re <= 1'd0;
    csrbank27_ev_enable0_we <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 3'd7))) begin
        csrbank27_ev_enable0_re <= interface27_bank_bus_we;
        csrbank27_ev_enable0_we <= csrbank27_re;
    end
end
assign csrbank27_clocks_per_tick0_r = interface27_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank27_clocks_per_tick0_we <= 1'd0;
    csrbank27_clocks_per_tick0_re <= 1'd0;
    if ((csrbank27_sel & (interface27_bank_bus_adr[9:0] == 4'd8))) begin
        csrbank27_clocks_per_tick0_re <= interface27_bank_bus_we;
        csrbank27_clocks_per_tick0_we <= csrbank27_re;
    end
end
always @(*) begin
    ticktimer_reset <= 1'd0;
    if (ticktimer_control_re) begin
        ticktimer_reset <= ticktimer_control_storage;
    end
end
assign csrbank27_control0_w = ticktimer_control_storage;
assign csrbank27_time1_w = ticktimer_time_status[63:32];
assign csrbank27_time0_w = ticktimer_time_status[31:0];
assign ticktimer_time_we = csrbank27_time0_we;
assign csrbank27_msleep_target1_w = ticktimer_msleep_target_storage[63:32];
assign csrbank27_msleep_target0_w = ticktimer_msleep_target_storage[31:0];
assign ticktimer_status_status = ticktimer_alarm0;
assign csrbank27_ev_status_w = ticktimer_status_status;
assign ticktimer_status_we = csrbank27_ev_status_we;
assign ticktimer_pending_status = ticktimer_alarm1;
assign csrbank27_ev_pending_w = ticktimer_pending_status;
assign ticktimer_pending_we = csrbank27_ev_pending_we;
assign ticktimer_alarm2 = ticktimer_enable_storage;
assign csrbank27_ev_enable0_w = ticktimer_enable_storage;
assign csrbank27_clocks_per_tick0_w = ticktimer_clocks_per_tick_storage[31:0];
assign csrbank28_sel = (interface28_bank_bus_adr[15:10] == 5'd28);
assign csrbank28_re = interface28_bank_bus_re;
assign csrbank28_load0_r = interface28_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank28_load0_re <= 1'd0;
    csrbank28_load0_we <= 1'd0;
    if ((csrbank28_sel & (interface28_bank_bus_adr[9:0] == 1'd0))) begin
        csrbank28_load0_re <= interface28_bank_bus_we;
        csrbank28_load0_we <= csrbank28_re;
    end
end
assign csrbank28_reload0_r = interface28_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank28_reload0_re <= 1'd0;
    csrbank28_reload0_we <= 1'd0;
    if ((csrbank28_sel & (interface28_bank_bus_adr[9:0] == 1'd1))) begin
        csrbank28_reload0_re <= interface28_bank_bus_we;
        csrbank28_reload0_we <= csrbank28_re;
    end
end
assign csrbank28_en0_r = interface28_bank_bus_dat_w[0];
always @(*) begin
    csrbank28_en0_we <= 1'd0;
    csrbank28_en0_re <= 1'd0;
    if ((csrbank28_sel & (interface28_bank_bus_adr[9:0] == 2'd2))) begin
        csrbank28_en0_re <= interface28_bank_bus_we;
        csrbank28_en0_we <= csrbank28_re;
    end
end
assign csrbank28_update_value0_r = interface28_bank_bus_dat_w[0];
always @(*) begin
    csrbank28_update_value0_re <= 1'd0;
    csrbank28_update_value0_we <= 1'd0;
    if ((csrbank28_sel & (interface28_bank_bus_adr[9:0] == 2'd3))) begin
        csrbank28_update_value0_re <= interface28_bank_bus_we;
        csrbank28_update_value0_we <= csrbank28_re;
    end
end
assign csrbank28_value_r = interface28_bank_bus_dat_w[31:0];
always @(*) begin
    csrbank28_value_we <= 1'd0;
    csrbank28_value_re <= 1'd0;
    if ((csrbank28_sel & (interface28_bank_bus_adr[9:0] == 3'd4))) begin
        csrbank28_value_re <= interface28_bank_bus_we;
        csrbank28_value_we <= csrbank28_re;
    end
end
assign csrbank28_ev_status_r = interface28_bank_bus_dat_w[0];
always @(*) begin
    csrbank28_ev_status_we <= 1'd0;
    csrbank28_ev_status_re <= 1'd0;
    if ((csrbank28_sel & (interface28_bank_bus_adr[9:0] == 3'd5))) begin
        csrbank28_ev_status_re <= interface28_bank_bus_we;
        csrbank28_ev_status_we <= csrbank28_re;
    end
end
assign csrbank28_ev_pending_r = interface28_bank_bus_dat_w[0];
always @(*) begin
    csrbank28_ev_pending_re <= 1'd0;
    csrbank28_ev_pending_we <= 1'd0;
    if ((csrbank28_sel & (interface28_bank_bus_adr[9:0] == 3'd6))) begin
        csrbank28_ev_pending_re <= interface28_bank_bus_we;
        csrbank28_ev_pending_we <= csrbank28_re;
    end
end
assign csrbank28_ev_enable0_r = interface28_bank_bus_dat_w[0];
always @(*) begin
    csrbank28_ev_enable0_re <= 1'd0;
    csrbank28_ev_enable0_we <= 1'd0;
    if ((csrbank28_sel & (interface28_bank_bus_adr[9:0] == 3'd7))) begin
        csrbank28_ev_enable0_re <= interface28_bank_bus_we;
        csrbank28_ev_enable0_we <= csrbank28_re;
    end
end
assign csrbank28_load0_w = cramsoc_load_storage[31:0];
assign csrbank28_reload0_w = cramsoc_reload_storage[31:0];
assign csrbank28_en0_w = cramsoc_en_storage;
assign csrbank28_update_value0_w = cramsoc_update_value_storage;
assign csrbank28_value_w = cramsoc_value_status[31:0];
assign cramsoc_value_we = csrbank28_value_we;
assign cramsoc_status_status = cramsoc_zero0;
assign csrbank28_ev_status_w = cramsoc_status_status;
assign cramsoc_status_we = csrbank28_ev_status_we;
assign cramsoc_pending_status = cramsoc_zero1;
assign csrbank28_ev_pending_w = cramsoc_pending_status;
assign cramsoc_pending_we = csrbank28_ev_pending_we;
assign cramsoc_zero2 = cramsoc_enable_storage;
assign csrbank28_ev_enable0_w = cramsoc_enable_storage;
assign csr_interconnect_adr = cramsoc_adr;
assign csr_interconnect_we = cramsoc_we;
assign csr_interconnect_dat_w = cramsoc_dat_w;
assign csr_interconnect_re = cramsoc_re;
assign cramsoc_dat_r = csr_interconnect_dat_r;
assign interface0_bank_bus_adr = csr_interconnect_adr;
assign interface1_bank_bus_adr = csr_interconnect_adr;
assign interface2_bank_bus_adr = csr_interconnect_adr;
assign interface3_bank_bus_adr = csr_interconnect_adr;
assign interface4_bank_bus_adr = csr_interconnect_adr;
assign interface5_bank_bus_adr = csr_interconnect_adr;
assign interface6_bank_bus_adr = csr_interconnect_adr;
assign interface7_bank_bus_adr = csr_interconnect_adr;
assign interface8_bank_bus_adr = csr_interconnect_adr;
assign interface9_bank_bus_adr = csr_interconnect_adr;
assign interface10_bank_bus_adr = csr_interconnect_adr;
assign interface11_bank_bus_adr = csr_interconnect_adr;
assign interface12_bank_bus_adr = csr_interconnect_adr;
assign interface13_bank_bus_adr = csr_interconnect_adr;
assign interface14_bank_bus_adr = csr_interconnect_adr;
assign interface15_bank_bus_adr = csr_interconnect_adr;
assign interface16_bank_bus_adr = csr_interconnect_adr;
assign interface17_bank_bus_adr = csr_interconnect_adr;
assign interface18_bank_bus_adr = csr_interconnect_adr;
assign interface19_bank_bus_adr = csr_interconnect_adr;
assign interface20_bank_bus_adr = csr_interconnect_adr;
assign interface21_bank_bus_adr = csr_interconnect_adr;
assign interface22_bank_bus_adr = csr_interconnect_adr;
assign interface23_bank_bus_adr = csr_interconnect_adr;
assign interface24_bank_bus_adr = csr_interconnect_adr;
assign interface25_bank_bus_adr = csr_interconnect_adr;
assign interface26_bank_bus_adr = csr_interconnect_adr;
assign interface27_bank_bus_adr = csr_interconnect_adr;
assign interface28_bank_bus_adr = csr_interconnect_adr;
assign interface0_bank_bus_we = csr_interconnect_we;
assign interface1_bank_bus_we = csr_interconnect_we;
assign interface2_bank_bus_we = csr_interconnect_we;
assign interface3_bank_bus_we = csr_interconnect_we;
assign interface4_bank_bus_we = csr_interconnect_we;
assign interface5_bank_bus_we = csr_interconnect_we;
assign interface6_bank_bus_we = csr_interconnect_we;
assign interface7_bank_bus_we = csr_interconnect_we;
assign interface8_bank_bus_we = csr_interconnect_we;
assign interface9_bank_bus_we = csr_interconnect_we;
assign interface10_bank_bus_we = csr_interconnect_we;
assign interface11_bank_bus_we = csr_interconnect_we;
assign interface12_bank_bus_we = csr_interconnect_we;
assign interface13_bank_bus_we = csr_interconnect_we;
assign interface14_bank_bus_we = csr_interconnect_we;
assign interface15_bank_bus_we = csr_interconnect_we;
assign interface16_bank_bus_we = csr_interconnect_we;
assign interface17_bank_bus_we = csr_interconnect_we;
assign interface18_bank_bus_we = csr_interconnect_we;
assign interface19_bank_bus_we = csr_interconnect_we;
assign interface20_bank_bus_we = csr_interconnect_we;
assign interface21_bank_bus_we = csr_interconnect_we;
assign interface22_bank_bus_we = csr_interconnect_we;
assign interface23_bank_bus_we = csr_interconnect_we;
assign interface24_bank_bus_we = csr_interconnect_we;
assign interface25_bank_bus_we = csr_interconnect_we;
assign interface26_bank_bus_we = csr_interconnect_we;
assign interface27_bank_bus_we = csr_interconnect_we;
assign interface28_bank_bus_we = csr_interconnect_we;
assign interface0_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface1_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface2_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface3_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface4_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface5_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface6_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface7_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface8_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface9_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface10_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface11_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface12_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface13_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface14_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface15_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface16_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface17_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface18_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface19_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface20_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface21_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface22_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface23_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface24_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface25_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface26_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface27_bank_bus_dat_w = csr_interconnect_dat_w;
assign interface28_bank_bus_dat_w = csr_interconnect_dat_w;
assign csr_interconnect_dat_r = ((((((((((((((((((((((((((((interface0_bank_bus_dat_r | interface1_bank_bus_dat_r) | interface2_bank_bus_dat_r) | interface3_bank_bus_dat_r) | interface4_bank_bus_dat_r) | interface5_bank_bus_dat_r) | interface6_bank_bus_dat_r) | interface7_bank_bus_dat_r) | interface8_bank_bus_dat_r) | interface9_bank_bus_dat_r) | interface10_bank_bus_dat_r) | interface11_bank_bus_dat_r) | interface12_bank_bus_dat_r) | interface13_bank_bus_dat_r) | interface14_bank_bus_dat_r) | interface15_bank_bus_dat_r) | interface16_bank_bus_dat_r) | interface17_bank_bus_dat_r) | interface18_bank_bus_dat_r) | interface19_bank_bus_dat_r) | interface20_bank_bus_dat_r) | interface21_bank_bus_dat_r) | interface22_bank_bus_dat_r) | interface23_bank_bus_dat_r) | interface24_bank_bus_dat_r) | interface25_bank_bus_dat_r) | interface26_bank_bus_dat_r) | interface27_bank_bus_dat_r) | interface28_bank_bus_dat_r);
assign interface0_bank_bus_re = csr_interconnect_re;
assign interface1_bank_bus_re = csr_interconnect_re;
assign interface2_bank_bus_re = csr_interconnect_re;
assign interface3_bank_bus_re = csr_interconnect_re;
assign interface4_bank_bus_re = csr_interconnect_re;
assign interface5_bank_bus_re = csr_interconnect_re;
assign interface6_bank_bus_re = csr_interconnect_re;
assign interface7_bank_bus_re = csr_interconnect_re;
assign interface8_bank_bus_re = csr_interconnect_re;
assign interface9_bank_bus_re = csr_interconnect_re;
assign interface10_bank_bus_re = csr_interconnect_re;
assign interface11_bank_bus_re = csr_interconnect_re;
assign interface12_bank_bus_re = csr_interconnect_re;
assign interface13_bank_bus_re = csr_interconnect_re;
assign interface14_bank_bus_re = csr_interconnect_re;
assign interface15_bank_bus_re = csr_interconnect_re;
assign interface16_bank_bus_re = csr_interconnect_re;
assign interface17_bank_bus_re = csr_interconnect_re;
assign interface18_bank_bus_re = csr_interconnect_re;
assign interface19_bank_bus_re = csr_interconnect_re;
assign interface20_bank_bus_re = csr_interconnect_re;
assign interface21_bank_bus_re = csr_interconnect_re;
assign interface22_bank_bus_re = csr_interconnect_re;
assign interface23_bank_bus_re = csr_interconnect_re;
assign interface24_bank_bus_re = csr_interconnect_re;
assign interface25_bank_bus_re = csr_interconnect_re;
assign interface26_bank_bus_re = csr_interconnect_re;
assign interface27_bank_bus_re = csr_interconnect_re;
assign interface28_bank_bus_re = csr_interconnect_re;
assign slice_proxy0 = cramsoc_corecsr_aw_payload_addr[31:2];
assign slice_proxy1 = cramsoc_corecsr_ar_payload_addr[31:2];
always @(*) begin
    array_muxed0 <= 1'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed0 <= socbushandler_aw_valid;
        end
    endcase
end
always @(*) begin
    array_muxed1 <= 1'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed1 <= socbushandler_aw_first;
        end
    endcase
end
always @(*) begin
    array_muxed2 <= 1'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed2 <= socbushandler_aw_last;
        end
    endcase
end
always @(*) begin
    array_muxed3 <= 32'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed3 <= socbushandler_aw_payload_addr;
        end
    endcase
end
always @(*) begin
    array_muxed4 <= 3'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed4 <= socbushandler_aw_payload_prot;
        end
    endcase
end
always @(*) begin
    array_muxed5 <= 1'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed5 <= socbushandler_w_valid;
        end
    endcase
end
always @(*) begin
    array_muxed6 <= 1'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed6 <= socbushandler_w_first;
        end
    endcase
end
always @(*) begin
    array_muxed7 <= 1'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed7 <= socbushandler_w_last;
        end
    endcase
end
always @(*) begin
    array_muxed8 <= 32'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed8 <= socbushandler_w_payload_data;
        end
    endcase
end
always @(*) begin
    array_muxed9 <= 4'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed9 <= socbushandler_w_payload_strb;
        end
    endcase
end
always @(*) begin
    array_muxed10 <= 1'd0;
    case (socbushandler_rr_write_grant)
        default: begin
            array_muxed10 <= socbushandler_b_ready;
        end
    endcase
end
always @(*) begin
    array_muxed11 <= 1'd0;
    case (socbushandler_rr_read_grant)
        default: begin
            array_muxed11 <= socbushandler_ar_valid;
        end
    endcase
end
always @(*) begin
    array_muxed12 <= 1'd0;
    case (socbushandler_rr_read_grant)
        default: begin
            array_muxed12 <= socbushandler_ar_first;
        end
    endcase
end
always @(*) begin
    array_muxed13 <= 1'd0;
    case (socbushandler_rr_read_grant)
        default: begin
            array_muxed13 <= socbushandler_ar_last;
        end
    endcase
end
always @(*) begin
    array_muxed14 <= 32'd0;
    case (socbushandler_rr_read_grant)
        default: begin
            array_muxed14 <= socbushandler_ar_payload_addr;
        end
    endcase
end
always @(*) begin
    array_muxed15 <= 3'd0;
    case (socbushandler_rr_read_grant)
        default: begin
            array_muxed15 <= socbushandler_ar_payload_prot;
        end
    endcase
end
always @(*) begin
    array_muxed16 <= 1'd0;
    case (socbushandler_rr_read_grant)
        default: begin
            array_muxed16 <= socbushandler_r_ready;
        end
    endcase
end
assign ticktimer_pause1 = multiregimpl0_regs1;
assign ticktimer_load_xfer_ps_toggle_o = multiregimpl1_regs1;
assign ticktimer_load_xfer_ps_ack_toggle_o = multiregimpl2_regs1;
assign ticktimer_paused0 = multiregimpl3_regs1;
assign ticktimer_timer_sync_ping_toggle_o = multiregimpl4_regs1;
assign ticktimer_timer_sync_pong_toggle_o = multiregimpl5_regs1;
assign ticktimer_timer_sync_obuffer = multiregimpl6_regs1;
assign ticktimer_resume_sync_ping_toggle_o = multiregimpl7_regs1;
assign ticktimer_resume_sync_pong_toggle_o = multiregimpl8_regs1;
assign ticktimer_resume_sync_obuffer = multiregimpl9_regs1;
assign ticktimer_reset_xfer_ps_toggle_o = multiregimpl10_regs1;
assign ticktimer_reset_xfer_ps_ack_toggle_o = multiregimpl11_regs1;
assign ticktimer_ping_ps_toggle_o = multiregimpl12_regs1;
assign ticktimer_ping_ps_ack_toggle_o = multiregimpl13_regs1;
assign ticktimer_pong_ps_toggle_o = multiregimpl14_regs1;
assign ticktimer_pong_ps_ack_toggle_o = multiregimpl15_regs1;
assign ticktimer_target_xfer_ping_toggle_o = multiregimpl16_regs1;
assign ticktimer_target_xfer_pong_toggle_o = multiregimpl17_regs1;
assign ticktimer_target_xfer_obuffer = multiregimpl18_regs1;


//------------------------------------------------------------------------------
// Synchronous Logic
//------------------------------------------------------------------------------

always @(posedge always_on_clk) begin
    cpu_int_active <= (cramsoc_interrupt == {1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0, 1'd0});
    irqarray0_eventsourceflex0_trigger_d <= irqarray0_interrupts[0];
    if ((irqarray0_eventsourceflex0_trigger_filtered | irqarray0_trigger[0])) begin
        irqarray0_eventsourceflex0_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex0_clear) begin
            irqarray0_eventsourceflex0_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex0_pending <= irqarray0_eventsourceflex0_pending;
        end
    end
    irqarray0_eventsourceflex1_trigger_d <= irqarray0_interrupts[1];
    if ((irqarray0_eventsourceflex1_trigger_filtered | irqarray0_trigger[1])) begin
        irqarray0_eventsourceflex1_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex1_clear) begin
            irqarray0_eventsourceflex1_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex1_pending <= irqarray0_eventsourceflex1_pending;
        end
    end
    irqarray0_eventsourceflex2_trigger_d <= irqarray0_interrupts[2];
    if ((irqarray0_eventsourceflex2_trigger_filtered | irqarray0_trigger[2])) begin
        irqarray0_eventsourceflex2_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex2_clear) begin
            irqarray0_eventsourceflex2_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex2_pending <= irqarray0_eventsourceflex2_pending;
        end
    end
    irqarray0_eventsourceflex3_trigger_d <= irqarray0_interrupts[3];
    if ((irqarray0_eventsourceflex3_trigger_filtered | irqarray0_trigger[3])) begin
        irqarray0_eventsourceflex3_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex3_clear) begin
            irqarray0_eventsourceflex3_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex3_pending <= irqarray0_eventsourceflex3_pending;
        end
    end
    irqarray0_eventsourceflex4_trigger_d <= irqarray0_interrupts[4];
    if ((irqarray0_eventsourceflex4_trigger_filtered | irqarray0_trigger[4])) begin
        irqarray0_eventsourceflex4_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex4_clear) begin
            irqarray0_eventsourceflex4_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex4_pending <= irqarray0_eventsourceflex4_pending;
        end
    end
    irqarray0_eventsourceflex5_trigger_d <= irqarray0_interrupts[5];
    if ((irqarray0_eventsourceflex5_trigger_filtered | irqarray0_trigger[5])) begin
        irqarray0_eventsourceflex5_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex5_clear) begin
            irqarray0_eventsourceflex5_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex5_pending <= irqarray0_eventsourceflex5_pending;
        end
    end
    irqarray0_eventsourceflex6_trigger_d <= irqarray0_interrupts[6];
    if ((irqarray0_eventsourceflex6_trigger_filtered | irqarray0_trigger[6])) begin
        irqarray0_eventsourceflex6_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex6_clear) begin
            irqarray0_eventsourceflex6_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex6_pending <= irqarray0_eventsourceflex6_pending;
        end
    end
    irqarray0_eventsourceflex7_trigger_d <= irqarray0_interrupts[7];
    if ((irqarray0_eventsourceflex7_trigger_filtered | irqarray0_trigger[7])) begin
        irqarray0_eventsourceflex7_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex7_clear) begin
            irqarray0_eventsourceflex7_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex7_pending <= irqarray0_eventsourceflex7_pending;
        end
    end
    irqarray0_eventsourceflex8_trigger_d <= irqarray0_interrupts[8];
    if ((irqarray0_eventsourceflex8_trigger_filtered | irqarray0_trigger[8])) begin
        irqarray0_eventsourceflex8_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex8_clear) begin
            irqarray0_eventsourceflex8_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex8_pending <= irqarray0_eventsourceflex8_pending;
        end
    end
    irqarray0_eventsourceflex9_trigger_d <= irqarray0_interrupts[9];
    if ((irqarray0_eventsourceflex9_trigger_filtered | irqarray0_trigger[9])) begin
        irqarray0_eventsourceflex9_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex9_clear) begin
            irqarray0_eventsourceflex9_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex9_pending <= irqarray0_eventsourceflex9_pending;
        end
    end
    irqarray0_eventsourceflex10_trigger_d <= irqarray0_interrupts[10];
    if ((irqarray0_eventsourceflex10_trigger_filtered | irqarray0_trigger[10])) begin
        irqarray0_eventsourceflex10_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex10_clear) begin
            irqarray0_eventsourceflex10_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex10_pending <= irqarray0_eventsourceflex10_pending;
        end
    end
    irqarray0_eventsourceflex11_trigger_d <= irqarray0_interrupts[11];
    if ((irqarray0_eventsourceflex11_trigger_filtered | irqarray0_trigger[11])) begin
        irqarray0_eventsourceflex11_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex11_clear) begin
            irqarray0_eventsourceflex11_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex11_pending <= irqarray0_eventsourceflex11_pending;
        end
    end
    irqarray0_eventsourceflex12_trigger_d <= irqarray0_interrupts[12];
    if ((irqarray0_eventsourceflex12_trigger_filtered | irqarray0_trigger[12])) begin
        irqarray0_eventsourceflex12_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex12_clear) begin
            irqarray0_eventsourceflex12_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex12_pending <= irqarray0_eventsourceflex12_pending;
        end
    end
    irqarray0_eventsourceflex13_trigger_d <= irqarray0_interrupts[13];
    if ((irqarray0_eventsourceflex13_trigger_filtered | irqarray0_trigger[13])) begin
        irqarray0_eventsourceflex13_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex13_clear) begin
            irqarray0_eventsourceflex13_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex13_pending <= irqarray0_eventsourceflex13_pending;
        end
    end
    irqarray0_eventsourceflex14_trigger_d <= irqarray0_interrupts[14];
    if ((irqarray0_eventsourceflex14_trigger_filtered | irqarray0_trigger[14])) begin
        irqarray0_eventsourceflex14_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex14_clear) begin
            irqarray0_eventsourceflex14_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex14_pending <= irqarray0_eventsourceflex14_pending;
        end
    end
    irqarray0_eventsourceflex15_trigger_d <= irqarray0_interrupts[15];
    if ((irqarray0_eventsourceflex15_trigger_filtered | irqarray0_trigger[15])) begin
        irqarray0_eventsourceflex15_pending <= 1'd1;
    end else begin
        if (irqarray0_eventsourceflex15_clear) begin
            irqarray0_eventsourceflex15_pending <= 1'd0;
        end else begin
            irqarray0_eventsourceflex15_pending <= irqarray0_eventsourceflex15_pending;
        end
    end
    irqarray1_eventsourceflex16_trigger_d <= irqarray1_interrupts[0];
    if ((irqarray1_eventsourceflex16_trigger_filtered | irqarray1_trigger[0])) begin
        irqarray1_eventsourceflex16_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex16_clear) begin
            irqarray1_eventsourceflex16_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex16_pending <= irqarray1_eventsourceflex16_pending;
        end
    end
    irqarray1_eventsourceflex17_trigger_d <= irqarray1_interrupts[1];
    if ((irqarray1_eventsourceflex17_trigger_filtered | irqarray1_trigger[1])) begin
        irqarray1_eventsourceflex17_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex17_clear) begin
            irqarray1_eventsourceflex17_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex17_pending <= irqarray1_eventsourceflex17_pending;
        end
    end
    irqarray1_eventsourceflex18_trigger_d <= irqarray1_interrupts[2];
    if ((irqarray1_eventsourceflex18_trigger_filtered | irqarray1_trigger[2])) begin
        irqarray1_eventsourceflex18_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex18_clear) begin
            irqarray1_eventsourceflex18_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex18_pending <= irqarray1_eventsourceflex18_pending;
        end
    end
    irqarray1_eventsourceflex19_trigger_d <= irqarray1_interrupts[3];
    if ((irqarray1_eventsourceflex19_trigger_filtered | irqarray1_trigger[3])) begin
        irqarray1_eventsourceflex19_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex19_clear) begin
            irqarray1_eventsourceflex19_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex19_pending <= irqarray1_eventsourceflex19_pending;
        end
    end
    irqarray1_eventsourceflex20_trigger_d <= irqarray1_interrupts[4];
    if ((irqarray1_eventsourceflex20_trigger_filtered | irqarray1_trigger[4])) begin
        irqarray1_eventsourceflex20_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex20_clear) begin
            irqarray1_eventsourceflex20_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex20_pending <= irqarray1_eventsourceflex20_pending;
        end
    end
    irqarray1_eventsourceflex21_trigger_d <= irqarray1_interrupts[5];
    if ((irqarray1_eventsourceflex21_trigger_filtered | irqarray1_trigger[5])) begin
        irqarray1_eventsourceflex21_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex21_clear) begin
            irqarray1_eventsourceflex21_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex21_pending <= irqarray1_eventsourceflex21_pending;
        end
    end
    irqarray1_eventsourceflex22_trigger_d <= irqarray1_interrupts[6];
    if ((irqarray1_eventsourceflex22_trigger_filtered | irqarray1_trigger[6])) begin
        irqarray1_eventsourceflex22_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex22_clear) begin
            irqarray1_eventsourceflex22_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex22_pending <= irqarray1_eventsourceflex22_pending;
        end
    end
    irqarray1_eventsourceflex23_trigger_d <= irqarray1_interrupts[7];
    if ((irqarray1_eventsourceflex23_trigger_filtered | irqarray1_trigger[7])) begin
        irqarray1_eventsourceflex23_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex23_clear) begin
            irqarray1_eventsourceflex23_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex23_pending <= irqarray1_eventsourceflex23_pending;
        end
    end
    irqarray1_eventsourceflex24_trigger_d <= irqarray1_interrupts[8];
    if ((irqarray1_eventsourceflex24_trigger_filtered | irqarray1_trigger[8])) begin
        irqarray1_eventsourceflex24_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex24_clear) begin
            irqarray1_eventsourceflex24_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex24_pending <= irqarray1_eventsourceflex24_pending;
        end
    end
    irqarray1_eventsourceflex25_trigger_d <= irqarray1_interrupts[9];
    if ((irqarray1_eventsourceflex25_trigger_filtered | irqarray1_trigger[9])) begin
        irqarray1_eventsourceflex25_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex25_clear) begin
            irqarray1_eventsourceflex25_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex25_pending <= irqarray1_eventsourceflex25_pending;
        end
    end
    irqarray1_eventsourceflex26_trigger_d <= irqarray1_interrupts[10];
    if ((irqarray1_eventsourceflex26_trigger_filtered | irqarray1_trigger[10])) begin
        irqarray1_eventsourceflex26_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex26_clear) begin
            irqarray1_eventsourceflex26_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex26_pending <= irqarray1_eventsourceflex26_pending;
        end
    end
    irqarray1_eventsourceflex27_trigger_d <= irqarray1_interrupts[11];
    if ((irqarray1_eventsourceflex27_trigger_filtered | irqarray1_trigger[11])) begin
        irqarray1_eventsourceflex27_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex27_clear) begin
            irqarray1_eventsourceflex27_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex27_pending <= irqarray1_eventsourceflex27_pending;
        end
    end
    irqarray1_eventsourceflex28_trigger_d <= irqarray1_interrupts[12];
    if ((irqarray1_eventsourceflex28_trigger_filtered | irqarray1_trigger[12])) begin
        irqarray1_eventsourceflex28_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex28_clear) begin
            irqarray1_eventsourceflex28_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex28_pending <= irqarray1_eventsourceflex28_pending;
        end
    end
    irqarray1_eventsourceflex29_trigger_d <= irqarray1_interrupts[13];
    if ((irqarray1_eventsourceflex29_trigger_filtered | irqarray1_trigger[13])) begin
        irqarray1_eventsourceflex29_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex29_clear) begin
            irqarray1_eventsourceflex29_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex29_pending <= irqarray1_eventsourceflex29_pending;
        end
    end
    irqarray1_eventsourceflex30_trigger_d <= irqarray1_interrupts[14];
    if ((irqarray1_eventsourceflex30_trigger_filtered | irqarray1_trigger[14])) begin
        irqarray1_eventsourceflex30_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex30_clear) begin
            irqarray1_eventsourceflex30_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex30_pending <= irqarray1_eventsourceflex30_pending;
        end
    end
    irqarray1_eventsourceflex31_trigger_d <= irqarray1_interrupts[15];
    if ((irqarray1_eventsourceflex31_trigger_filtered | irqarray1_trigger[15])) begin
        irqarray1_eventsourceflex31_pending <= 1'd1;
    end else begin
        if (irqarray1_eventsourceflex31_clear) begin
            irqarray1_eventsourceflex31_pending <= 1'd0;
        end else begin
            irqarray1_eventsourceflex31_pending <= irqarray1_eventsourceflex31_pending;
        end
    end
    irqarray2_eventsourceflex32_trigger_d <= irqarray2_interrupts[0];
    if ((irqarray2_eventsourceflex32_trigger_filtered | irqarray2_trigger[0])) begin
        irqarray2_eventsourceflex32_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex32_clear) begin
            irqarray2_eventsourceflex32_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex32_pending <= irqarray2_eventsourceflex32_pending;
        end
    end
    irqarray2_eventsourceflex33_trigger_d <= irqarray2_interrupts[1];
    if ((irqarray2_eventsourceflex33_trigger_filtered | irqarray2_trigger[1])) begin
        irqarray2_eventsourceflex33_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex33_clear) begin
            irqarray2_eventsourceflex33_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex33_pending <= irqarray2_eventsourceflex33_pending;
        end
    end
    irqarray2_eventsourceflex34_trigger_d <= irqarray2_interrupts[2];
    if ((irqarray2_eventsourceflex34_trigger_filtered | irqarray2_trigger[2])) begin
        irqarray2_eventsourceflex34_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex34_clear) begin
            irqarray2_eventsourceflex34_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex34_pending <= irqarray2_eventsourceflex34_pending;
        end
    end
    irqarray2_eventsourceflex35_trigger_d <= irqarray2_interrupts[3];
    if ((irqarray2_eventsourceflex35_trigger_filtered | irqarray2_trigger[3])) begin
        irqarray2_eventsourceflex35_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex35_clear) begin
            irqarray2_eventsourceflex35_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex35_pending <= irqarray2_eventsourceflex35_pending;
        end
    end
    irqarray2_eventsourceflex36_trigger_d <= irqarray2_interrupts[4];
    if ((irqarray2_eventsourceflex36_trigger_filtered | irqarray2_trigger[4])) begin
        irqarray2_eventsourceflex36_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex36_clear) begin
            irqarray2_eventsourceflex36_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex36_pending <= irqarray2_eventsourceflex36_pending;
        end
    end
    irqarray2_eventsourceflex37_trigger_d <= irqarray2_interrupts[5];
    if ((irqarray2_eventsourceflex37_trigger_filtered | irqarray2_trigger[5])) begin
        irqarray2_eventsourceflex37_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex37_clear) begin
            irqarray2_eventsourceflex37_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex37_pending <= irqarray2_eventsourceflex37_pending;
        end
    end
    irqarray2_eventsourceflex38_trigger_d <= irqarray2_interrupts[6];
    if ((irqarray2_eventsourceflex38_trigger_filtered | irqarray2_trigger[6])) begin
        irqarray2_eventsourceflex38_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex38_clear) begin
            irqarray2_eventsourceflex38_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex38_pending <= irqarray2_eventsourceflex38_pending;
        end
    end
    irqarray2_eventsourceflex39_trigger_d <= irqarray2_interrupts[7];
    if ((irqarray2_eventsourceflex39_trigger_filtered | irqarray2_trigger[7])) begin
        irqarray2_eventsourceflex39_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex39_clear) begin
            irqarray2_eventsourceflex39_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex39_pending <= irqarray2_eventsourceflex39_pending;
        end
    end
    irqarray2_eventsourceflex40_trigger_d <= irqarray2_interrupts[8];
    if ((irqarray2_eventsourceflex40_trigger_filtered | irqarray2_trigger[8])) begin
        irqarray2_eventsourceflex40_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex40_clear) begin
            irqarray2_eventsourceflex40_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex40_pending <= irqarray2_eventsourceflex40_pending;
        end
    end
    irqarray2_eventsourceflex41_trigger_d <= irqarray2_interrupts[9];
    if ((irqarray2_eventsourceflex41_trigger_filtered | irqarray2_trigger[9])) begin
        irqarray2_eventsourceflex41_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex41_clear) begin
            irqarray2_eventsourceflex41_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex41_pending <= irqarray2_eventsourceflex41_pending;
        end
    end
    irqarray2_eventsourceflex42_trigger_d <= irqarray2_interrupts[10];
    if ((irqarray2_eventsourceflex42_trigger_filtered | irqarray2_trigger[10])) begin
        irqarray2_eventsourceflex42_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex42_clear) begin
            irqarray2_eventsourceflex42_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex42_pending <= irqarray2_eventsourceflex42_pending;
        end
    end
    irqarray2_eventsourceflex43_trigger_d <= irqarray2_interrupts[11];
    if ((irqarray2_eventsourceflex43_trigger_filtered | irqarray2_trigger[11])) begin
        irqarray2_eventsourceflex43_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex43_clear) begin
            irqarray2_eventsourceflex43_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex43_pending <= irqarray2_eventsourceflex43_pending;
        end
    end
    irqarray2_eventsourceflex44_trigger_d <= irqarray2_interrupts[12];
    if ((irqarray2_eventsourceflex44_trigger_filtered | irqarray2_trigger[12])) begin
        irqarray2_eventsourceflex44_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex44_clear) begin
            irqarray2_eventsourceflex44_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex44_pending <= irqarray2_eventsourceflex44_pending;
        end
    end
    irqarray2_eventsourceflex45_trigger_d <= irqarray2_interrupts[13];
    if ((irqarray2_eventsourceflex45_trigger_filtered | irqarray2_trigger[13])) begin
        irqarray2_eventsourceflex45_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex45_clear) begin
            irqarray2_eventsourceflex45_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex45_pending <= irqarray2_eventsourceflex45_pending;
        end
    end
    irqarray2_eventsourceflex46_trigger_d <= irqarray2_interrupts[14];
    if ((irqarray2_eventsourceflex46_trigger_filtered | irqarray2_trigger[14])) begin
        irqarray2_eventsourceflex46_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex46_clear) begin
            irqarray2_eventsourceflex46_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex46_pending <= irqarray2_eventsourceflex46_pending;
        end
    end
    irqarray2_eventsourceflex47_trigger_d <= irqarray2_interrupts[15];
    if ((irqarray2_eventsourceflex47_trigger_filtered | irqarray2_trigger[15])) begin
        irqarray2_eventsourceflex47_pending <= 1'd1;
    end else begin
        if (irqarray2_eventsourceflex47_clear) begin
            irqarray2_eventsourceflex47_pending <= 1'd0;
        end else begin
            irqarray2_eventsourceflex47_pending <= irqarray2_eventsourceflex47_pending;
        end
    end
    irqarray3_eventsourceflex48_trigger_d <= irqarray3_interrupts[0];
    if ((irqarray3_eventsourceflex48_trigger_filtered | irqarray3_trigger[0])) begin
        irqarray3_eventsourceflex48_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex48_clear) begin
            irqarray3_eventsourceflex48_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex48_pending <= irqarray3_eventsourceflex48_pending;
        end
    end
    irqarray3_eventsourceflex49_trigger_d <= irqarray3_interrupts[1];
    if ((irqarray3_eventsourceflex49_trigger_filtered | irqarray3_trigger[1])) begin
        irqarray3_eventsourceflex49_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex49_clear) begin
            irqarray3_eventsourceflex49_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex49_pending <= irqarray3_eventsourceflex49_pending;
        end
    end
    irqarray3_eventsourceflex50_trigger_d <= irqarray3_interrupts[2];
    if ((irqarray3_eventsourceflex50_trigger_filtered | irqarray3_trigger[2])) begin
        irqarray3_eventsourceflex50_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex50_clear) begin
            irqarray3_eventsourceflex50_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex50_pending <= irqarray3_eventsourceflex50_pending;
        end
    end
    irqarray3_eventsourceflex51_trigger_d <= irqarray3_interrupts[3];
    if ((irqarray3_eventsourceflex51_trigger_filtered | irqarray3_trigger[3])) begin
        irqarray3_eventsourceflex51_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex51_clear) begin
            irqarray3_eventsourceflex51_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex51_pending <= irqarray3_eventsourceflex51_pending;
        end
    end
    irqarray3_eventsourceflex52_trigger_d <= irqarray3_interrupts[4];
    if ((irqarray3_eventsourceflex52_trigger_filtered | irqarray3_trigger[4])) begin
        irqarray3_eventsourceflex52_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex52_clear) begin
            irqarray3_eventsourceflex52_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex52_pending <= irqarray3_eventsourceflex52_pending;
        end
    end
    irqarray3_eventsourceflex53_trigger_d <= irqarray3_interrupts[5];
    if ((irqarray3_eventsourceflex53_trigger_filtered | irqarray3_trigger[5])) begin
        irqarray3_eventsourceflex53_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex53_clear) begin
            irqarray3_eventsourceflex53_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex53_pending <= irqarray3_eventsourceflex53_pending;
        end
    end
    irqarray3_eventsourceflex54_trigger_d <= irqarray3_interrupts[6];
    if ((irqarray3_eventsourceflex54_trigger_filtered | irqarray3_trigger[6])) begin
        irqarray3_eventsourceflex54_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex54_clear) begin
            irqarray3_eventsourceflex54_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex54_pending <= irqarray3_eventsourceflex54_pending;
        end
    end
    irqarray3_eventsourceflex55_trigger_d <= irqarray3_interrupts[7];
    if ((irqarray3_eventsourceflex55_trigger_filtered | irqarray3_trigger[7])) begin
        irqarray3_eventsourceflex55_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex55_clear) begin
            irqarray3_eventsourceflex55_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex55_pending <= irqarray3_eventsourceflex55_pending;
        end
    end
    irqarray3_eventsourceflex56_trigger_d <= irqarray3_interrupts[8];
    if ((irqarray3_eventsourceflex56_trigger_filtered | irqarray3_trigger[8])) begin
        irqarray3_eventsourceflex56_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex56_clear) begin
            irqarray3_eventsourceflex56_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex56_pending <= irqarray3_eventsourceflex56_pending;
        end
    end
    irqarray3_eventsourceflex57_trigger_d <= irqarray3_interrupts[9];
    if ((irqarray3_eventsourceflex57_trigger_filtered | irqarray3_trigger[9])) begin
        irqarray3_eventsourceflex57_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex57_clear) begin
            irqarray3_eventsourceflex57_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex57_pending <= irqarray3_eventsourceflex57_pending;
        end
    end
    irqarray3_eventsourceflex58_trigger_d <= irqarray3_interrupts[10];
    if ((irqarray3_eventsourceflex58_trigger_filtered | irqarray3_trigger[10])) begin
        irqarray3_eventsourceflex58_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex58_clear) begin
            irqarray3_eventsourceflex58_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex58_pending <= irqarray3_eventsourceflex58_pending;
        end
    end
    irqarray3_eventsourceflex59_trigger_d <= irqarray3_interrupts[11];
    if ((irqarray3_eventsourceflex59_trigger_filtered | irqarray3_trigger[11])) begin
        irqarray3_eventsourceflex59_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex59_clear) begin
            irqarray3_eventsourceflex59_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex59_pending <= irqarray3_eventsourceflex59_pending;
        end
    end
    irqarray3_eventsourceflex60_trigger_d <= irqarray3_interrupts[12];
    if ((irqarray3_eventsourceflex60_trigger_filtered | irqarray3_trigger[12])) begin
        irqarray3_eventsourceflex60_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex60_clear) begin
            irqarray3_eventsourceflex60_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex60_pending <= irqarray3_eventsourceflex60_pending;
        end
    end
    irqarray3_eventsourceflex61_trigger_d <= irqarray3_interrupts[13];
    if ((irqarray3_eventsourceflex61_trigger_filtered | irqarray3_trigger[13])) begin
        irqarray3_eventsourceflex61_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex61_clear) begin
            irqarray3_eventsourceflex61_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex61_pending <= irqarray3_eventsourceflex61_pending;
        end
    end
    irqarray3_eventsourceflex62_trigger_d <= irqarray3_interrupts[14];
    if ((irqarray3_eventsourceflex62_trigger_filtered | irqarray3_trigger[14])) begin
        irqarray3_eventsourceflex62_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex62_clear) begin
            irqarray3_eventsourceflex62_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex62_pending <= irqarray3_eventsourceflex62_pending;
        end
    end
    irqarray3_eventsourceflex63_trigger_d <= irqarray3_interrupts[15];
    if ((irqarray3_eventsourceflex63_trigger_filtered | irqarray3_trigger[15])) begin
        irqarray3_eventsourceflex63_pending <= 1'd1;
    end else begin
        if (irqarray3_eventsourceflex63_clear) begin
            irqarray3_eventsourceflex63_pending <= 1'd0;
        end else begin
            irqarray3_eventsourceflex63_pending <= irqarray3_eventsourceflex63_pending;
        end
    end
    irqarray4_eventsourceflex64_trigger_d <= irqarray4_interrupts[0];
    if ((irqarray4_eventsourceflex64_trigger_filtered | irqarray4_trigger[0])) begin
        irqarray4_eventsourceflex64_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex64_clear) begin
            irqarray4_eventsourceflex64_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex64_pending <= irqarray4_eventsourceflex64_pending;
        end
    end
    irqarray4_eventsourceflex65_trigger_d <= irqarray4_interrupts[1];
    if ((irqarray4_eventsourceflex65_trigger_filtered | irqarray4_trigger[1])) begin
        irqarray4_eventsourceflex65_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex65_clear) begin
            irqarray4_eventsourceflex65_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex65_pending <= irqarray4_eventsourceflex65_pending;
        end
    end
    irqarray4_eventsourceflex66_trigger_d <= irqarray4_interrupts[2];
    if ((irqarray4_eventsourceflex66_trigger_filtered | irqarray4_trigger[2])) begin
        irqarray4_eventsourceflex66_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex66_clear) begin
            irqarray4_eventsourceflex66_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex66_pending <= irqarray4_eventsourceflex66_pending;
        end
    end
    irqarray4_eventsourceflex67_trigger_d <= irqarray4_interrupts[3];
    if ((irqarray4_eventsourceflex67_trigger_filtered | irqarray4_trigger[3])) begin
        irqarray4_eventsourceflex67_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex67_clear) begin
            irqarray4_eventsourceflex67_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex67_pending <= irqarray4_eventsourceflex67_pending;
        end
    end
    irqarray4_eventsourceflex68_trigger_d <= irqarray4_interrupts[4];
    if ((irqarray4_eventsourceflex68_trigger_filtered | irqarray4_trigger[4])) begin
        irqarray4_eventsourceflex68_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex68_clear) begin
            irqarray4_eventsourceflex68_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex68_pending <= irqarray4_eventsourceflex68_pending;
        end
    end
    irqarray4_eventsourceflex69_trigger_d <= irqarray4_interrupts[5];
    if ((irqarray4_eventsourceflex69_trigger_filtered | irqarray4_trigger[5])) begin
        irqarray4_eventsourceflex69_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex69_clear) begin
            irqarray4_eventsourceflex69_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex69_pending <= irqarray4_eventsourceflex69_pending;
        end
    end
    irqarray4_eventsourceflex70_trigger_d <= irqarray4_interrupts[6];
    if ((irqarray4_eventsourceflex70_trigger_filtered | irqarray4_trigger[6])) begin
        irqarray4_eventsourceflex70_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex70_clear) begin
            irqarray4_eventsourceflex70_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex70_pending <= irqarray4_eventsourceflex70_pending;
        end
    end
    irqarray4_eventsourceflex71_trigger_d <= irqarray4_interrupts[7];
    if ((irqarray4_eventsourceflex71_trigger_filtered | irqarray4_trigger[7])) begin
        irqarray4_eventsourceflex71_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex71_clear) begin
            irqarray4_eventsourceflex71_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex71_pending <= irqarray4_eventsourceflex71_pending;
        end
    end
    irqarray4_eventsourceflex72_trigger_d <= irqarray4_interrupts[8];
    if ((irqarray4_eventsourceflex72_trigger_filtered | irqarray4_trigger[8])) begin
        irqarray4_eventsourceflex72_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex72_clear) begin
            irqarray4_eventsourceflex72_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex72_pending <= irqarray4_eventsourceflex72_pending;
        end
    end
    irqarray4_eventsourceflex73_trigger_d <= irqarray4_interrupts[9];
    if ((irqarray4_eventsourceflex73_trigger_filtered | irqarray4_trigger[9])) begin
        irqarray4_eventsourceflex73_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex73_clear) begin
            irqarray4_eventsourceflex73_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex73_pending <= irqarray4_eventsourceflex73_pending;
        end
    end
    irqarray4_eventsourceflex74_trigger_d <= irqarray4_interrupts[10];
    if ((irqarray4_eventsourceflex74_trigger_filtered | irqarray4_trigger[10])) begin
        irqarray4_eventsourceflex74_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex74_clear) begin
            irqarray4_eventsourceflex74_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex74_pending <= irqarray4_eventsourceflex74_pending;
        end
    end
    irqarray4_eventsourceflex75_trigger_d <= irqarray4_interrupts[11];
    if ((irqarray4_eventsourceflex75_trigger_filtered | irqarray4_trigger[11])) begin
        irqarray4_eventsourceflex75_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex75_clear) begin
            irqarray4_eventsourceflex75_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex75_pending <= irqarray4_eventsourceflex75_pending;
        end
    end
    irqarray4_eventsourceflex76_trigger_d <= irqarray4_interrupts[12];
    if ((irqarray4_eventsourceflex76_trigger_filtered | irqarray4_trigger[12])) begin
        irqarray4_eventsourceflex76_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex76_clear) begin
            irqarray4_eventsourceflex76_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex76_pending <= irqarray4_eventsourceflex76_pending;
        end
    end
    irqarray4_eventsourceflex77_trigger_d <= irqarray4_interrupts[13];
    if ((irqarray4_eventsourceflex77_trigger_filtered | irqarray4_trigger[13])) begin
        irqarray4_eventsourceflex77_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex77_clear) begin
            irqarray4_eventsourceflex77_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex77_pending <= irqarray4_eventsourceflex77_pending;
        end
    end
    irqarray4_eventsourceflex78_trigger_d <= irqarray4_interrupts[14];
    if ((irqarray4_eventsourceflex78_trigger_filtered | irqarray4_trigger[14])) begin
        irqarray4_eventsourceflex78_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex78_clear) begin
            irqarray4_eventsourceflex78_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex78_pending <= irqarray4_eventsourceflex78_pending;
        end
    end
    irqarray4_eventsourceflex79_trigger_d <= irqarray4_interrupts[15];
    if ((irqarray4_eventsourceflex79_trigger_filtered | irqarray4_trigger[15])) begin
        irqarray4_eventsourceflex79_pending <= 1'd1;
    end else begin
        if (irqarray4_eventsourceflex79_clear) begin
            irqarray4_eventsourceflex79_pending <= 1'd0;
        end else begin
            irqarray4_eventsourceflex79_pending <= irqarray4_eventsourceflex79_pending;
        end
    end
    irqarray5_eventsourceflex80_trigger_d <= irqarray5_interrupts[0];
    if ((irqarray5_eventsourceflex80_trigger_filtered | irqarray5_trigger[0])) begin
        irqarray5_eventsourceflex80_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex80_clear) begin
            irqarray5_eventsourceflex80_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex80_pending <= irqarray5_eventsourceflex80_pending;
        end
    end
    irqarray5_eventsourceflex81_trigger_d <= irqarray5_interrupts[1];
    if ((irqarray5_eventsourceflex81_trigger_filtered | irqarray5_trigger[1])) begin
        irqarray5_eventsourceflex81_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex81_clear) begin
            irqarray5_eventsourceflex81_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex81_pending <= irqarray5_eventsourceflex81_pending;
        end
    end
    irqarray5_eventsourceflex82_trigger_d <= irqarray5_interrupts[2];
    if ((irqarray5_eventsourceflex82_trigger_filtered | irqarray5_trigger[2])) begin
        irqarray5_eventsourceflex82_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex82_clear) begin
            irqarray5_eventsourceflex82_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex82_pending <= irqarray5_eventsourceflex82_pending;
        end
    end
    irqarray5_eventsourceflex83_trigger_d <= irqarray5_interrupts[3];
    if ((irqarray5_eventsourceflex83_trigger_filtered | irqarray5_trigger[3])) begin
        irqarray5_eventsourceflex83_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex83_clear) begin
            irqarray5_eventsourceflex83_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex83_pending <= irqarray5_eventsourceflex83_pending;
        end
    end
    irqarray5_eventsourceflex84_trigger_d <= irqarray5_interrupts[4];
    if ((irqarray5_eventsourceflex84_trigger_filtered | irqarray5_trigger[4])) begin
        irqarray5_eventsourceflex84_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex84_clear) begin
            irqarray5_eventsourceflex84_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex84_pending <= irqarray5_eventsourceflex84_pending;
        end
    end
    irqarray5_eventsourceflex85_trigger_d <= irqarray5_interrupts[5];
    if ((irqarray5_eventsourceflex85_trigger_filtered | irqarray5_trigger[5])) begin
        irqarray5_eventsourceflex85_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex85_clear) begin
            irqarray5_eventsourceflex85_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex85_pending <= irqarray5_eventsourceflex85_pending;
        end
    end
    irqarray5_eventsourceflex86_trigger_d <= irqarray5_interrupts[6];
    if ((irqarray5_eventsourceflex86_trigger_filtered | irqarray5_trigger[6])) begin
        irqarray5_eventsourceflex86_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex86_clear) begin
            irqarray5_eventsourceflex86_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex86_pending <= irqarray5_eventsourceflex86_pending;
        end
    end
    irqarray5_eventsourceflex87_trigger_d <= irqarray5_interrupts[7];
    if ((irqarray5_eventsourceflex87_trigger_filtered | irqarray5_trigger[7])) begin
        irqarray5_eventsourceflex87_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex87_clear) begin
            irqarray5_eventsourceflex87_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex87_pending <= irqarray5_eventsourceflex87_pending;
        end
    end
    irqarray5_eventsourceflex88_trigger_d <= irqarray5_interrupts[8];
    if ((irqarray5_eventsourceflex88_trigger_filtered | irqarray5_trigger[8])) begin
        irqarray5_eventsourceflex88_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex88_clear) begin
            irqarray5_eventsourceflex88_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex88_pending <= irqarray5_eventsourceflex88_pending;
        end
    end
    irqarray5_eventsourceflex89_trigger_d <= irqarray5_interrupts[9];
    if ((irqarray5_eventsourceflex89_trigger_filtered | irqarray5_trigger[9])) begin
        irqarray5_eventsourceflex89_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex89_clear) begin
            irqarray5_eventsourceflex89_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex89_pending <= irqarray5_eventsourceflex89_pending;
        end
    end
    irqarray5_eventsourceflex90_trigger_d <= irqarray5_interrupts[10];
    if ((irqarray5_eventsourceflex90_trigger_filtered | irqarray5_trigger[10])) begin
        irqarray5_eventsourceflex90_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex90_clear) begin
            irqarray5_eventsourceflex90_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex90_pending <= irqarray5_eventsourceflex90_pending;
        end
    end
    irqarray5_eventsourceflex91_trigger_d <= irqarray5_interrupts[11];
    if ((irqarray5_eventsourceflex91_trigger_filtered | irqarray5_trigger[11])) begin
        irqarray5_eventsourceflex91_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex91_clear) begin
            irqarray5_eventsourceflex91_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex91_pending <= irqarray5_eventsourceflex91_pending;
        end
    end
    irqarray5_eventsourceflex92_trigger_d <= irqarray5_interrupts[12];
    if ((irqarray5_eventsourceflex92_trigger_filtered | irqarray5_trigger[12])) begin
        irqarray5_eventsourceflex92_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex92_clear) begin
            irqarray5_eventsourceflex92_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex92_pending <= irqarray5_eventsourceflex92_pending;
        end
    end
    irqarray5_eventsourceflex93_trigger_d <= irqarray5_interrupts[13];
    if ((irqarray5_eventsourceflex93_trigger_filtered | irqarray5_trigger[13])) begin
        irqarray5_eventsourceflex93_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex93_clear) begin
            irqarray5_eventsourceflex93_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex93_pending <= irqarray5_eventsourceflex93_pending;
        end
    end
    irqarray5_eventsourceflex94_trigger_d <= irqarray5_interrupts[14];
    if ((irqarray5_eventsourceflex94_trigger_filtered | irqarray5_trigger[14])) begin
        irqarray5_eventsourceflex94_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex94_clear) begin
            irqarray5_eventsourceflex94_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex94_pending <= irqarray5_eventsourceflex94_pending;
        end
    end
    irqarray5_eventsourceflex95_trigger_d <= irqarray5_interrupts[15];
    if ((irqarray5_eventsourceflex95_trigger_filtered | irqarray5_trigger[15])) begin
        irqarray5_eventsourceflex95_pending <= 1'd1;
    end else begin
        if (irqarray5_eventsourceflex95_clear) begin
            irqarray5_eventsourceflex95_pending <= 1'd0;
        end else begin
            irqarray5_eventsourceflex95_pending <= irqarray5_eventsourceflex95_pending;
        end
    end
    irqarray6_eventsourceflex96_trigger_d <= irqarray6_interrupts[0];
    if ((irqarray6_eventsourceflex96_trigger_filtered | irqarray6_trigger[0])) begin
        irqarray6_eventsourceflex96_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex96_clear) begin
            irqarray6_eventsourceflex96_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex96_pending <= irqarray6_eventsourceflex96_pending;
        end
    end
    irqarray6_eventsourceflex97_trigger_d <= irqarray6_interrupts[1];
    if ((irqarray6_eventsourceflex97_trigger_filtered | irqarray6_trigger[1])) begin
        irqarray6_eventsourceflex97_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex97_clear) begin
            irqarray6_eventsourceflex97_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex97_pending <= irqarray6_eventsourceflex97_pending;
        end
    end
    irqarray6_eventsourceflex98_trigger_d <= irqarray6_interrupts[2];
    if ((irqarray6_eventsourceflex98_trigger_filtered | irqarray6_trigger[2])) begin
        irqarray6_eventsourceflex98_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex98_clear) begin
            irqarray6_eventsourceflex98_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex98_pending <= irqarray6_eventsourceflex98_pending;
        end
    end
    irqarray6_eventsourceflex99_trigger_d <= irqarray6_interrupts[3];
    if ((irqarray6_eventsourceflex99_trigger_filtered | irqarray6_trigger[3])) begin
        irqarray6_eventsourceflex99_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex99_clear) begin
            irqarray6_eventsourceflex99_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex99_pending <= irqarray6_eventsourceflex99_pending;
        end
    end
    irqarray6_eventsourceflex100_trigger_d <= irqarray6_interrupts[4];
    if ((irqarray6_eventsourceflex100_trigger_filtered | irqarray6_trigger[4])) begin
        irqarray6_eventsourceflex100_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex100_clear) begin
            irqarray6_eventsourceflex100_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex100_pending <= irqarray6_eventsourceflex100_pending;
        end
    end
    irqarray6_eventsourceflex101_trigger_d <= irqarray6_interrupts[5];
    if ((irqarray6_eventsourceflex101_trigger_filtered | irqarray6_trigger[5])) begin
        irqarray6_eventsourceflex101_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex101_clear) begin
            irqarray6_eventsourceflex101_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex101_pending <= irqarray6_eventsourceflex101_pending;
        end
    end
    irqarray6_eventsourceflex102_trigger_d <= irqarray6_interrupts[6];
    if ((irqarray6_eventsourceflex102_trigger_filtered | irqarray6_trigger[6])) begin
        irqarray6_eventsourceflex102_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex102_clear) begin
            irqarray6_eventsourceflex102_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex102_pending <= irqarray6_eventsourceflex102_pending;
        end
    end
    irqarray6_eventsourceflex103_trigger_d <= irqarray6_interrupts[7];
    if ((irqarray6_eventsourceflex103_trigger_filtered | irqarray6_trigger[7])) begin
        irqarray6_eventsourceflex103_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex103_clear) begin
            irqarray6_eventsourceflex103_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex103_pending <= irqarray6_eventsourceflex103_pending;
        end
    end
    irqarray6_eventsourceflex104_trigger_d <= irqarray6_interrupts[8];
    if ((irqarray6_eventsourceflex104_trigger_filtered | irqarray6_trigger[8])) begin
        irqarray6_eventsourceflex104_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex104_clear) begin
            irqarray6_eventsourceflex104_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex104_pending <= irqarray6_eventsourceflex104_pending;
        end
    end
    irqarray6_eventsourceflex105_trigger_d <= irqarray6_interrupts[9];
    if ((irqarray6_eventsourceflex105_trigger_filtered | irqarray6_trigger[9])) begin
        irqarray6_eventsourceflex105_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex105_clear) begin
            irqarray6_eventsourceflex105_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex105_pending <= irqarray6_eventsourceflex105_pending;
        end
    end
    irqarray6_eventsourceflex106_trigger_d <= irqarray6_interrupts[10];
    if ((irqarray6_eventsourceflex106_trigger_filtered | irqarray6_trigger[10])) begin
        irqarray6_eventsourceflex106_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex106_clear) begin
            irqarray6_eventsourceflex106_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex106_pending <= irqarray6_eventsourceflex106_pending;
        end
    end
    irqarray6_eventsourceflex107_trigger_d <= irqarray6_interrupts[11];
    if ((irqarray6_eventsourceflex107_trigger_filtered | irqarray6_trigger[11])) begin
        irqarray6_eventsourceflex107_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex107_clear) begin
            irqarray6_eventsourceflex107_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex107_pending <= irqarray6_eventsourceflex107_pending;
        end
    end
    irqarray6_eventsourceflex108_trigger_d <= irqarray6_interrupts[12];
    if ((irqarray6_eventsourceflex108_trigger_filtered | irqarray6_trigger[12])) begin
        irqarray6_eventsourceflex108_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex108_clear) begin
            irqarray6_eventsourceflex108_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex108_pending <= irqarray6_eventsourceflex108_pending;
        end
    end
    irqarray6_eventsourceflex109_trigger_d <= irqarray6_interrupts[13];
    if ((irqarray6_eventsourceflex109_trigger_filtered | irqarray6_trigger[13])) begin
        irqarray6_eventsourceflex109_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex109_clear) begin
            irqarray6_eventsourceflex109_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex109_pending <= irqarray6_eventsourceflex109_pending;
        end
    end
    irqarray6_eventsourceflex110_trigger_d <= irqarray6_interrupts[14];
    if ((irqarray6_eventsourceflex110_trigger_filtered | irqarray6_trigger[14])) begin
        irqarray6_eventsourceflex110_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex110_clear) begin
            irqarray6_eventsourceflex110_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex110_pending <= irqarray6_eventsourceflex110_pending;
        end
    end
    irqarray6_eventsourceflex111_trigger_d <= irqarray6_interrupts[15];
    if ((irqarray6_eventsourceflex111_trigger_filtered | irqarray6_trigger[15])) begin
        irqarray6_eventsourceflex111_pending <= 1'd1;
    end else begin
        if (irqarray6_eventsourceflex111_clear) begin
            irqarray6_eventsourceflex111_pending <= 1'd0;
        end else begin
            irqarray6_eventsourceflex111_pending <= irqarray6_eventsourceflex111_pending;
        end
    end
    irqarray7_eventsourceflex112_trigger_d <= irqarray7_interrupts[0];
    if ((irqarray7_eventsourceflex112_trigger_filtered | irqarray7_trigger[0])) begin
        irqarray7_eventsourceflex112_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex112_clear) begin
            irqarray7_eventsourceflex112_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex112_pending <= irqarray7_eventsourceflex112_pending;
        end
    end
    irqarray7_eventsourceflex113_trigger_d <= irqarray7_interrupts[1];
    if ((irqarray7_eventsourceflex113_trigger_filtered | irqarray7_trigger[1])) begin
        irqarray7_eventsourceflex113_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex113_clear) begin
            irqarray7_eventsourceflex113_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex113_pending <= irqarray7_eventsourceflex113_pending;
        end
    end
    irqarray7_eventsourceflex114_trigger_d <= irqarray7_interrupts[2];
    if ((irqarray7_eventsourceflex114_trigger_filtered | irqarray7_trigger[2])) begin
        irqarray7_eventsourceflex114_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex114_clear) begin
            irqarray7_eventsourceflex114_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex114_pending <= irqarray7_eventsourceflex114_pending;
        end
    end
    irqarray7_eventsourceflex115_trigger_d <= irqarray7_interrupts[3];
    if ((irqarray7_eventsourceflex115_trigger_filtered | irqarray7_trigger[3])) begin
        irqarray7_eventsourceflex115_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex115_clear) begin
            irqarray7_eventsourceflex115_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex115_pending <= irqarray7_eventsourceflex115_pending;
        end
    end
    irqarray7_eventsourceflex116_trigger_d <= irqarray7_interrupts[4];
    if ((irqarray7_eventsourceflex116_trigger_filtered | irqarray7_trigger[4])) begin
        irqarray7_eventsourceflex116_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex116_clear) begin
            irqarray7_eventsourceflex116_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex116_pending <= irqarray7_eventsourceflex116_pending;
        end
    end
    irqarray7_eventsourceflex117_trigger_d <= irqarray7_interrupts[5];
    if ((irqarray7_eventsourceflex117_trigger_filtered | irqarray7_trigger[5])) begin
        irqarray7_eventsourceflex117_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex117_clear) begin
            irqarray7_eventsourceflex117_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex117_pending <= irqarray7_eventsourceflex117_pending;
        end
    end
    irqarray7_eventsourceflex118_trigger_d <= irqarray7_interrupts[6];
    if ((irqarray7_eventsourceflex118_trigger_filtered | irqarray7_trigger[6])) begin
        irqarray7_eventsourceflex118_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex118_clear) begin
            irqarray7_eventsourceflex118_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex118_pending <= irqarray7_eventsourceflex118_pending;
        end
    end
    irqarray7_eventsourceflex119_trigger_d <= irqarray7_interrupts[7];
    if ((irqarray7_eventsourceflex119_trigger_filtered | irqarray7_trigger[7])) begin
        irqarray7_eventsourceflex119_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex119_clear) begin
            irqarray7_eventsourceflex119_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex119_pending <= irqarray7_eventsourceflex119_pending;
        end
    end
    irqarray7_eventsourceflex120_trigger_d <= irqarray7_interrupts[8];
    if ((irqarray7_eventsourceflex120_trigger_filtered | irqarray7_trigger[8])) begin
        irqarray7_eventsourceflex120_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex120_clear) begin
            irqarray7_eventsourceflex120_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex120_pending <= irqarray7_eventsourceflex120_pending;
        end
    end
    irqarray7_eventsourceflex121_trigger_d <= irqarray7_interrupts[9];
    if ((irqarray7_eventsourceflex121_trigger_filtered | irqarray7_trigger[9])) begin
        irqarray7_eventsourceflex121_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex121_clear) begin
            irqarray7_eventsourceflex121_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex121_pending <= irqarray7_eventsourceflex121_pending;
        end
    end
    irqarray7_eventsourceflex122_trigger_d <= irqarray7_interrupts[10];
    if ((irqarray7_eventsourceflex122_trigger_filtered | irqarray7_trigger[10])) begin
        irqarray7_eventsourceflex122_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex122_clear) begin
            irqarray7_eventsourceflex122_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex122_pending <= irqarray7_eventsourceflex122_pending;
        end
    end
    irqarray7_eventsourceflex123_trigger_d <= irqarray7_interrupts[11];
    if ((irqarray7_eventsourceflex123_trigger_filtered | irqarray7_trigger[11])) begin
        irqarray7_eventsourceflex123_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex123_clear) begin
            irqarray7_eventsourceflex123_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex123_pending <= irqarray7_eventsourceflex123_pending;
        end
    end
    irqarray7_eventsourceflex124_trigger_d <= irqarray7_interrupts[12];
    if ((irqarray7_eventsourceflex124_trigger_filtered | irqarray7_trigger[12])) begin
        irqarray7_eventsourceflex124_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex124_clear) begin
            irqarray7_eventsourceflex124_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex124_pending <= irqarray7_eventsourceflex124_pending;
        end
    end
    irqarray7_eventsourceflex125_trigger_d <= irqarray7_interrupts[13];
    if ((irqarray7_eventsourceflex125_trigger_filtered | irqarray7_trigger[13])) begin
        irqarray7_eventsourceflex125_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex125_clear) begin
            irqarray7_eventsourceflex125_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex125_pending <= irqarray7_eventsourceflex125_pending;
        end
    end
    irqarray7_eventsourceflex126_trigger_d <= irqarray7_interrupts[14];
    if ((irqarray7_eventsourceflex126_trigger_filtered | irqarray7_trigger[14])) begin
        irqarray7_eventsourceflex126_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex126_clear) begin
            irqarray7_eventsourceflex126_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex126_pending <= irqarray7_eventsourceflex126_pending;
        end
    end
    irqarray7_eventsourceflex127_trigger_d <= irqarray7_interrupts[15];
    if ((irqarray7_eventsourceflex127_trigger_filtered | irqarray7_trigger[15])) begin
        irqarray7_eventsourceflex127_pending <= 1'd1;
    end else begin
        if (irqarray7_eventsourceflex127_clear) begin
            irqarray7_eventsourceflex127_pending <= 1'd0;
        end else begin
            irqarray7_eventsourceflex127_pending <= irqarray7_eventsourceflex127_pending;
        end
    end
    irqarray8_eventsourceflex128_trigger_d <= irqarray8_interrupts[0];
    if ((irqarray8_eventsourceflex128_trigger_filtered | irqarray8_trigger[0])) begin
        irqarray8_eventsourceflex128_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex128_clear) begin
            irqarray8_eventsourceflex128_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex128_pending <= irqarray8_eventsourceflex128_pending;
        end
    end
    irqarray8_eventsourceflex129_trigger_d <= irqarray8_interrupts[1];
    if ((irqarray8_eventsourceflex129_trigger_filtered | irqarray8_trigger[1])) begin
        irqarray8_eventsourceflex129_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex129_clear) begin
            irqarray8_eventsourceflex129_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex129_pending <= irqarray8_eventsourceflex129_pending;
        end
    end
    irqarray8_eventsourceflex130_trigger_d <= irqarray8_interrupts[2];
    if ((irqarray8_eventsourceflex130_trigger_filtered | irqarray8_trigger[2])) begin
        irqarray8_eventsourceflex130_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex130_clear) begin
            irqarray8_eventsourceflex130_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex130_pending <= irqarray8_eventsourceflex130_pending;
        end
    end
    irqarray8_eventsourceflex131_trigger_d <= irqarray8_interrupts[3];
    if ((irqarray8_eventsourceflex131_trigger_filtered | irqarray8_trigger[3])) begin
        irqarray8_eventsourceflex131_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex131_clear) begin
            irqarray8_eventsourceflex131_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex131_pending <= irqarray8_eventsourceflex131_pending;
        end
    end
    irqarray8_eventsourceflex132_trigger_d <= irqarray8_interrupts[4];
    if ((irqarray8_eventsourceflex132_trigger_filtered | irqarray8_trigger[4])) begin
        irqarray8_eventsourceflex132_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex132_clear) begin
            irqarray8_eventsourceflex132_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex132_pending <= irqarray8_eventsourceflex132_pending;
        end
    end
    irqarray8_eventsourceflex133_trigger_d <= irqarray8_interrupts[5];
    if ((irqarray8_eventsourceflex133_trigger_filtered | irqarray8_trigger[5])) begin
        irqarray8_eventsourceflex133_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex133_clear) begin
            irqarray8_eventsourceflex133_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex133_pending <= irqarray8_eventsourceflex133_pending;
        end
    end
    irqarray8_eventsourceflex134_trigger_d <= irqarray8_interrupts[6];
    if ((irqarray8_eventsourceflex134_trigger_filtered | irqarray8_trigger[6])) begin
        irqarray8_eventsourceflex134_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex134_clear) begin
            irqarray8_eventsourceflex134_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex134_pending <= irqarray8_eventsourceflex134_pending;
        end
    end
    irqarray8_eventsourceflex135_trigger_d <= irqarray8_interrupts[7];
    if ((irqarray8_eventsourceflex135_trigger_filtered | irqarray8_trigger[7])) begin
        irqarray8_eventsourceflex135_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex135_clear) begin
            irqarray8_eventsourceflex135_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex135_pending <= irqarray8_eventsourceflex135_pending;
        end
    end
    irqarray8_eventsourceflex136_trigger_d <= irqarray8_interrupts[8];
    if ((irqarray8_eventsourceflex136_trigger_filtered | irqarray8_trigger[8])) begin
        irqarray8_eventsourceflex136_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex136_clear) begin
            irqarray8_eventsourceflex136_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex136_pending <= irqarray8_eventsourceflex136_pending;
        end
    end
    irqarray8_eventsourceflex137_trigger_d <= irqarray8_interrupts[9];
    if ((irqarray8_eventsourceflex137_trigger_filtered | irqarray8_trigger[9])) begin
        irqarray8_eventsourceflex137_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex137_clear) begin
            irqarray8_eventsourceflex137_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex137_pending <= irqarray8_eventsourceflex137_pending;
        end
    end
    irqarray8_eventsourceflex138_trigger_d <= irqarray8_interrupts[10];
    if ((irqarray8_eventsourceflex138_trigger_filtered | irqarray8_trigger[10])) begin
        irqarray8_eventsourceflex138_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex138_clear) begin
            irqarray8_eventsourceflex138_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex138_pending <= irqarray8_eventsourceflex138_pending;
        end
    end
    irqarray8_eventsourceflex139_trigger_d <= irqarray8_interrupts[11];
    if ((irqarray8_eventsourceflex139_trigger_filtered | irqarray8_trigger[11])) begin
        irqarray8_eventsourceflex139_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex139_clear) begin
            irqarray8_eventsourceflex139_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex139_pending <= irqarray8_eventsourceflex139_pending;
        end
    end
    irqarray8_eventsourceflex140_trigger_d <= irqarray8_interrupts[12];
    if ((irqarray8_eventsourceflex140_trigger_filtered | irqarray8_trigger[12])) begin
        irqarray8_eventsourceflex140_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex140_clear) begin
            irqarray8_eventsourceflex140_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex140_pending <= irqarray8_eventsourceflex140_pending;
        end
    end
    irqarray8_eventsourceflex141_trigger_d <= irqarray8_interrupts[13];
    if ((irqarray8_eventsourceflex141_trigger_filtered | irqarray8_trigger[13])) begin
        irqarray8_eventsourceflex141_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex141_clear) begin
            irqarray8_eventsourceflex141_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex141_pending <= irqarray8_eventsourceflex141_pending;
        end
    end
    irqarray8_eventsourceflex142_trigger_d <= irqarray8_interrupts[14];
    if ((irqarray8_eventsourceflex142_trigger_filtered | irqarray8_trigger[14])) begin
        irqarray8_eventsourceflex142_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex142_clear) begin
            irqarray8_eventsourceflex142_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex142_pending <= irqarray8_eventsourceflex142_pending;
        end
    end
    irqarray8_eventsourceflex143_trigger_d <= irqarray8_interrupts[15];
    if ((irqarray8_eventsourceflex143_trigger_filtered | irqarray8_trigger[15])) begin
        irqarray8_eventsourceflex143_pending <= 1'd1;
    end else begin
        if (irqarray8_eventsourceflex143_clear) begin
            irqarray8_eventsourceflex143_pending <= 1'd0;
        end else begin
            irqarray8_eventsourceflex143_pending <= irqarray8_eventsourceflex143_pending;
        end
    end
    irqarray9_eventsourceflex144_trigger_d <= irqarray9_interrupts[0];
    if ((irqarray9_eventsourceflex144_trigger_filtered | irqarray9_trigger[0])) begin
        irqarray9_eventsourceflex144_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex144_clear) begin
            irqarray9_eventsourceflex144_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex144_pending <= irqarray9_eventsourceflex144_pending;
        end
    end
    irqarray9_eventsourceflex145_trigger_d <= irqarray9_interrupts[1];
    if ((irqarray9_eventsourceflex145_trigger_filtered | irqarray9_trigger[1])) begin
        irqarray9_eventsourceflex145_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex145_clear) begin
            irqarray9_eventsourceflex145_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex145_pending <= irqarray9_eventsourceflex145_pending;
        end
    end
    irqarray9_eventsourceflex146_trigger_d <= irqarray9_interrupts[2];
    if ((irqarray9_eventsourceflex146_trigger_filtered | irqarray9_trigger[2])) begin
        irqarray9_eventsourceflex146_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex146_clear) begin
            irqarray9_eventsourceflex146_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex146_pending <= irqarray9_eventsourceflex146_pending;
        end
    end
    irqarray9_eventsourceflex147_trigger_d <= irqarray9_interrupts[3];
    if ((irqarray9_eventsourceflex147_trigger_filtered | irqarray9_trigger[3])) begin
        irqarray9_eventsourceflex147_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex147_clear) begin
            irqarray9_eventsourceflex147_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex147_pending <= irqarray9_eventsourceflex147_pending;
        end
    end
    irqarray9_eventsourceflex148_trigger_d <= irqarray9_interrupts[4];
    if ((irqarray9_eventsourceflex148_trigger_filtered | irqarray9_trigger[4])) begin
        irqarray9_eventsourceflex148_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex148_clear) begin
            irqarray9_eventsourceflex148_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex148_pending <= irqarray9_eventsourceflex148_pending;
        end
    end
    irqarray9_eventsourceflex149_trigger_d <= irqarray9_interrupts[5];
    if ((irqarray9_eventsourceflex149_trigger_filtered | irqarray9_trigger[5])) begin
        irqarray9_eventsourceflex149_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex149_clear) begin
            irqarray9_eventsourceflex149_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex149_pending <= irqarray9_eventsourceflex149_pending;
        end
    end
    irqarray9_eventsourceflex150_trigger_d <= irqarray9_interrupts[6];
    if ((irqarray9_eventsourceflex150_trigger_filtered | irqarray9_trigger[6])) begin
        irqarray9_eventsourceflex150_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex150_clear) begin
            irqarray9_eventsourceflex150_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex150_pending <= irqarray9_eventsourceflex150_pending;
        end
    end
    irqarray9_eventsourceflex151_trigger_d <= irqarray9_interrupts[7];
    if ((irqarray9_eventsourceflex151_trigger_filtered | irqarray9_trigger[7])) begin
        irqarray9_eventsourceflex151_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex151_clear) begin
            irqarray9_eventsourceflex151_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex151_pending <= irqarray9_eventsourceflex151_pending;
        end
    end
    irqarray9_eventsourceflex152_trigger_d <= irqarray9_interrupts[8];
    if ((irqarray9_eventsourceflex152_trigger_filtered | irqarray9_trigger[8])) begin
        irqarray9_eventsourceflex152_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex152_clear) begin
            irqarray9_eventsourceflex152_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex152_pending <= irqarray9_eventsourceflex152_pending;
        end
    end
    irqarray9_eventsourceflex153_trigger_d <= irqarray9_interrupts[9];
    if ((irqarray9_eventsourceflex153_trigger_filtered | irqarray9_trigger[9])) begin
        irqarray9_eventsourceflex153_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex153_clear) begin
            irqarray9_eventsourceflex153_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex153_pending <= irqarray9_eventsourceflex153_pending;
        end
    end
    irqarray9_eventsourceflex154_trigger_d <= irqarray9_interrupts[10];
    if ((irqarray9_eventsourceflex154_trigger_filtered | irqarray9_trigger[10])) begin
        irqarray9_eventsourceflex154_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex154_clear) begin
            irqarray9_eventsourceflex154_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex154_pending <= irqarray9_eventsourceflex154_pending;
        end
    end
    irqarray9_eventsourceflex155_trigger_d <= irqarray9_interrupts[11];
    if ((irqarray9_eventsourceflex155_trigger_filtered | irqarray9_trigger[11])) begin
        irqarray9_eventsourceflex155_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex155_clear) begin
            irqarray9_eventsourceflex155_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex155_pending <= irqarray9_eventsourceflex155_pending;
        end
    end
    irqarray9_eventsourceflex156_trigger_d <= irqarray9_interrupts[12];
    if ((irqarray9_eventsourceflex156_trigger_filtered | irqarray9_trigger[12])) begin
        irqarray9_eventsourceflex156_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex156_clear) begin
            irqarray9_eventsourceflex156_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex156_pending <= irqarray9_eventsourceflex156_pending;
        end
    end
    irqarray9_eventsourceflex157_trigger_d <= irqarray9_interrupts[13];
    if ((irqarray9_eventsourceflex157_trigger_filtered | irqarray9_trigger[13])) begin
        irqarray9_eventsourceflex157_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex157_clear) begin
            irqarray9_eventsourceflex157_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex157_pending <= irqarray9_eventsourceflex157_pending;
        end
    end
    irqarray9_eventsourceflex158_trigger_d <= irqarray9_interrupts[14];
    if ((irqarray9_eventsourceflex158_trigger_filtered | irqarray9_trigger[14])) begin
        irqarray9_eventsourceflex158_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex158_clear) begin
            irqarray9_eventsourceflex158_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex158_pending <= irqarray9_eventsourceflex158_pending;
        end
    end
    irqarray9_eventsourceflex159_trigger_d <= irqarray9_interrupts[15];
    if ((irqarray9_eventsourceflex159_trigger_filtered | irqarray9_trigger[15])) begin
        irqarray9_eventsourceflex159_pending <= 1'd1;
    end else begin
        if (irqarray9_eventsourceflex159_clear) begin
            irqarray9_eventsourceflex159_pending <= 1'd0;
        end else begin
            irqarray9_eventsourceflex159_pending <= irqarray9_eventsourceflex159_pending;
        end
    end
    irqarray10_eventsourceflex160_trigger_d <= irqarray10_interrupts[0];
    if ((irqarray10_eventsourceflex160_trigger_filtered | irqarray10_trigger[0])) begin
        irqarray10_eventsourceflex160_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex160_clear) begin
            irqarray10_eventsourceflex160_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex160_pending <= irqarray10_eventsourceflex160_pending;
        end
    end
    irqarray10_eventsourceflex161_trigger_d <= irqarray10_interrupts[1];
    if ((irqarray10_eventsourceflex161_trigger_filtered | irqarray10_trigger[1])) begin
        irqarray10_eventsourceflex161_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex161_clear) begin
            irqarray10_eventsourceflex161_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex161_pending <= irqarray10_eventsourceflex161_pending;
        end
    end
    irqarray10_eventsourceflex162_trigger_d <= irqarray10_interrupts[2];
    if ((irqarray10_eventsourceflex162_trigger_filtered | irqarray10_trigger[2])) begin
        irqarray10_eventsourceflex162_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex162_clear) begin
            irqarray10_eventsourceflex162_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex162_pending <= irqarray10_eventsourceflex162_pending;
        end
    end
    irqarray10_eventsourceflex163_trigger_d <= irqarray10_interrupts[3];
    if ((irqarray10_eventsourceflex163_trigger_filtered | irqarray10_trigger[3])) begin
        irqarray10_eventsourceflex163_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex163_clear) begin
            irqarray10_eventsourceflex163_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex163_pending <= irqarray10_eventsourceflex163_pending;
        end
    end
    irqarray10_eventsourceflex164_trigger_d <= irqarray10_interrupts[4];
    if ((irqarray10_eventsourceflex164_trigger_filtered | irqarray10_trigger[4])) begin
        irqarray10_eventsourceflex164_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex164_clear) begin
            irqarray10_eventsourceflex164_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex164_pending <= irqarray10_eventsourceflex164_pending;
        end
    end
    irqarray10_eventsourceflex165_trigger_d <= irqarray10_interrupts[5];
    if ((irqarray10_eventsourceflex165_trigger_filtered | irqarray10_trigger[5])) begin
        irqarray10_eventsourceflex165_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex165_clear) begin
            irqarray10_eventsourceflex165_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex165_pending <= irqarray10_eventsourceflex165_pending;
        end
    end
    irqarray10_eventsourceflex166_trigger_d <= irqarray10_interrupts[6];
    if ((irqarray10_eventsourceflex166_trigger_filtered | irqarray10_trigger[6])) begin
        irqarray10_eventsourceflex166_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex166_clear) begin
            irqarray10_eventsourceflex166_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex166_pending <= irqarray10_eventsourceflex166_pending;
        end
    end
    irqarray10_eventsourceflex167_trigger_d <= irqarray10_interrupts[7];
    if ((irqarray10_eventsourceflex167_trigger_filtered | irqarray10_trigger[7])) begin
        irqarray10_eventsourceflex167_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex167_clear) begin
            irqarray10_eventsourceflex167_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex167_pending <= irqarray10_eventsourceflex167_pending;
        end
    end
    irqarray10_eventsourceflex168_trigger_d <= irqarray10_interrupts[8];
    if ((irqarray10_eventsourceflex168_trigger_filtered | irqarray10_trigger[8])) begin
        irqarray10_eventsourceflex168_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex168_clear) begin
            irqarray10_eventsourceflex168_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex168_pending <= irqarray10_eventsourceflex168_pending;
        end
    end
    irqarray10_eventsourceflex169_trigger_d <= irqarray10_interrupts[9];
    if ((irqarray10_eventsourceflex169_trigger_filtered | irqarray10_trigger[9])) begin
        irqarray10_eventsourceflex169_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex169_clear) begin
            irqarray10_eventsourceflex169_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex169_pending <= irqarray10_eventsourceflex169_pending;
        end
    end
    irqarray10_eventsourceflex170_trigger_d <= irqarray10_interrupts[10];
    if ((irqarray10_eventsourceflex170_trigger_filtered | irqarray10_trigger[10])) begin
        irqarray10_eventsourceflex170_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex170_clear) begin
            irqarray10_eventsourceflex170_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex170_pending <= irqarray10_eventsourceflex170_pending;
        end
    end
    irqarray10_eventsourceflex171_trigger_d <= irqarray10_interrupts[11];
    if ((irqarray10_eventsourceflex171_trigger_filtered | irqarray10_trigger[11])) begin
        irqarray10_eventsourceflex171_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex171_clear) begin
            irqarray10_eventsourceflex171_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex171_pending <= irqarray10_eventsourceflex171_pending;
        end
    end
    irqarray10_eventsourceflex172_trigger_d <= irqarray10_interrupts[12];
    if ((irqarray10_eventsourceflex172_trigger_filtered | irqarray10_trigger[12])) begin
        irqarray10_eventsourceflex172_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex172_clear) begin
            irqarray10_eventsourceflex172_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex172_pending <= irqarray10_eventsourceflex172_pending;
        end
    end
    irqarray10_eventsourceflex173_trigger_d <= irqarray10_interrupts[13];
    if ((irqarray10_eventsourceflex173_trigger_filtered | irqarray10_trigger[13])) begin
        irqarray10_eventsourceflex173_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex173_clear) begin
            irqarray10_eventsourceflex173_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex173_pending <= irqarray10_eventsourceflex173_pending;
        end
    end
    irqarray10_eventsourceflex174_trigger_d <= irqarray10_interrupts[14];
    if ((irqarray10_eventsourceflex174_trigger_filtered | irqarray10_trigger[14])) begin
        irqarray10_eventsourceflex174_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex174_clear) begin
            irqarray10_eventsourceflex174_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex174_pending <= irqarray10_eventsourceflex174_pending;
        end
    end
    irqarray10_eventsourceflex175_trigger_d <= irqarray10_interrupts[15];
    if ((irqarray10_eventsourceflex175_trigger_filtered | irqarray10_trigger[15])) begin
        irqarray10_eventsourceflex175_pending <= 1'd1;
    end else begin
        if (irqarray10_eventsourceflex175_clear) begin
            irqarray10_eventsourceflex175_pending <= 1'd0;
        end else begin
            irqarray10_eventsourceflex175_pending <= irqarray10_eventsourceflex175_pending;
        end
    end
    irqarray11_eventsourceflex176_trigger_d <= irqarray11_interrupts[0];
    if ((irqarray11_eventsourceflex176_trigger_filtered | irqarray11_trigger[0])) begin
        irqarray11_eventsourceflex176_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex176_clear) begin
            irqarray11_eventsourceflex176_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex176_pending <= irqarray11_eventsourceflex176_pending;
        end
    end
    irqarray11_eventsourceflex177_trigger_d <= irqarray11_interrupts[1];
    if ((irqarray11_eventsourceflex177_trigger_filtered | irqarray11_trigger[1])) begin
        irqarray11_eventsourceflex177_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex177_clear) begin
            irqarray11_eventsourceflex177_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex177_pending <= irqarray11_eventsourceflex177_pending;
        end
    end
    irqarray11_eventsourceflex178_trigger_d <= irqarray11_interrupts[2];
    if ((irqarray11_eventsourceflex178_trigger_filtered | irqarray11_trigger[2])) begin
        irqarray11_eventsourceflex178_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex178_clear) begin
            irqarray11_eventsourceflex178_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex178_pending <= irqarray11_eventsourceflex178_pending;
        end
    end
    irqarray11_eventsourceflex179_trigger_d <= irqarray11_interrupts[3];
    if ((irqarray11_eventsourceflex179_trigger_filtered | irqarray11_trigger[3])) begin
        irqarray11_eventsourceflex179_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex179_clear) begin
            irqarray11_eventsourceflex179_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex179_pending <= irqarray11_eventsourceflex179_pending;
        end
    end
    irqarray11_eventsourceflex180_trigger_d <= irqarray11_interrupts[4];
    if ((irqarray11_eventsourceflex180_trigger_filtered | irqarray11_trigger[4])) begin
        irqarray11_eventsourceflex180_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex180_clear) begin
            irqarray11_eventsourceflex180_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex180_pending <= irqarray11_eventsourceflex180_pending;
        end
    end
    irqarray11_eventsourceflex181_trigger_d <= irqarray11_interrupts[5];
    if ((irqarray11_eventsourceflex181_trigger_filtered | irqarray11_trigger[5])) begin
        irqarray11_eventsourceflex181_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex181_clear) begin
            irqarray11_eventsourceflex181_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex181_pending <= irqarray11_eventsourceflex181_pending;
        end
    end
    irqarray11_eventsourceflex182_trigger_d <= irqarray11_interrupts[6];
    if ((irqarray11_eventsourceflex182_trigger_filtered | irqarray11_trigger[6])) begin
        irqarray11_eventsourceflex182_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex182_clear) begin
            irqarray11_eventsourceflex182_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex182_pending <= irqarray11_eventsourceflex182_pending;
        end
    end
    irqarray11_eventsourceflex183_trigger_d <= irqarray11_interrupts[7];
    if ((irqarray11_eventsourceflex183_trigger_filtered | irqarray11_trigger[7])) begin
        irqarray11_eventsourceflex183_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex183_clear) begin
            irqarray11_eventsourceflex183_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex183_pending <= irqarray11_eventsourceflex183_pending;
        end
    end
    irqarray11_eventsourceflex184_trigger_d <= irqarray11_interrupts[8];
    if ((irqarray11_eventsourceflex184_trigger_filtered | irqarray11_trigger[8])) begin
        irqarray11_eventsourceflex184_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex184_clear) begin
            irqarray11_eventsourceflex184_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex184_pending <= irqarray11_eventsourceflex184_pending;
        end
    end
    irqarray11_eventsourceflex185_trigger_d <= irqarray11_interrupts[9];
    if ((irqarray11_eventsourceflex185_trigger_filtered | irqarray11_trigger[9])) begin
        irqarray11_eventsourceflex185_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex185_clear) begin
            irqarray11_eventsourceflex185_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex185_pending <= irqarray11_eventsourceflex185_pending;
        end
    end
    irqarray11_eventsourceflex186_trigger_d <= irqarray11_interrupts[10];
    if ((irqarray11_eventsourceflex186_trigger_filtered | irqarray11_trigger[10])) begin
        irqarray11_eventsourceflex186_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex186_clear) begin
            irqarray11_eventsourceflex186_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex186_pending <= irqarray11_eventsourceflex186_pending;
        end
    end
    irqarray11_eventsourceflex187_trigger_d <= irqarray11_interrupts[11];
    if ((irqarray11_eventsourceflex187_trigger_filtered | irqarray11_trigger[11])) begin
        irqarray11_eventsourceflex187_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex187_clear) begin
            irqarray11_eventsourceflex187_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex187_pending <= irqarray11_eventsourceflex187_pending;
        end
    end
    irqarray11_eventsourceflex188_trigger_d <= irqarray11_interrupts[12];
    if ((irqarray11_eventsourceflex188_trigger_filtered | irqarray11_trigger[12])) begin
        irqarray11_eventsourceflex188_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex188_clear) begin
            irqarray11_eventsourceflex188_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex188_pending <= irqarray11_eventsourceflex188_pending;
        end
    end
    irqarray11_eventsourceflex189_trigger_d <= irqarray11_interrupts[13];
    if ((irqarray11_eventsourceflex189_trigger_filtered | irqarray11_trigger[13])) begin
        irqarray11_eventsourceflex189_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex189_clear) begin
            irqarray11_eventsourceflex189_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex189_pending <= irqarray11_eventsourceflex189_pending;
        end
    end
    irqarray11_eventsourceflex190_trigger_d <= irqarray11_interrupts[14];
    if ((irqarray11_eventsourceflex190_trigger_filtered | irqarray11_trigger[14])) begin
        irqarray11_eventsourceflex190_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex190_clear) begin
            irqarray11_eventsourceflex190_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex190_pending <= irqarray11_eventsourceflex190_pending;
        end
    end
    irqarray11_eventsourceflex191_trigger_d <= irqarray11_interrupts[15];
    if ((irqarray11_eventsourceflex191_trigger_filtered | irqarray11_trigger[15])) begin
        irqarray11_eventsourceflex191_pending <= 1'd1;
    end else begin
        if (irqarray11_eventsourceflex191_clear) begin
            irqarray11_eventsourceflex191_pending <= 1'd0;
        end else begin
            irqarray11_eventsourceflex191_pending <= irqarray11_eventsourceflex191_pending;
        end
    end
    irqarray12_eventsourceflex192_trigger_d <= irqarray12_interrupts[0];
    if ((irqarray12_eventsourceflex192_trigger_filtered | irqarray12_trigger[0])) begin
        irqarray12_eventsourceflex192_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex192_clear) begin
            irqarray12_eventsourceflex192_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex192_pending <= irqarray12_eventsourceflex192_pending;
        end
    end
    irqarray12_eventsourceflex193_trigger_d <= irqarray12_interrupts[1];
    if ((irqarray12_eventsourceflex193_trigger_filtered | irqarray12_trigger[1])) begin
        irqarray12_eventsourceflex193_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex193_clear) begin
            irqarray12_eventsourceflex193_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex193_pending <= irqarray12_eventsourceflex193_pending;
        end
    end
    irqarray12_eventsourceflex194_trigger_d <= irqarray12_interrupts[2];
    if ((irqarray12_eventsourceflex194_trigger_filtered | irqarray12_trigger[2])) begin
        irqarray12_eventsourceflex194_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex194_clear) begin
            irqarray12_eventsourceflex194_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex194_pending <= irqarray12_eventsourceflex194_pending;
        end
    end
    irqarray12_eventsourceflex195_trigger_d <= irqarray12_interrupts[3];
    if ((irqarray12_eventsourceflex195_trigger_filtered | irqarray12_trigger[3])) begin
        irqarray12_eventsourceflex195_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex195_clear) begin
            irqarray12_eventsourceflex195_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex195_pending <= irqarray12_eventsourceflex195_pending;
        end
    end
    irqarray12_eventsourceflex196_trigger_d <= irqarray12_interrupts[4];
    if ((irqarray12_eventsourceflex196_trigger_filtered | irqarray12_trigger[4])) begin
        irqarray12_eventsourceflex196_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex196_clear) begin
            irqarray12_eventsourceflex196_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex196_pending <= irqarray12_eventsourceflex196_pending;
        end
    end
    irqarray12_eventsourceflex197_trigger_d <= irqarray12_interrupts[5];
    if ((irqarray12_eventsourceflex197_trigger_filtered | irqarray12_trigger[5])) begin
        irqarray12_eventsourceflex197_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex197_clear) begin
            irqarray12_eventsourceflex197_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex197_pending <= irqarray12_eventsourceflex197_pending;
        end
    end
    irqarray12_eventsourceflex198_trigger_d <= irqarray12_interrupts[6];
    if ((irqarray12_eventsourceflex198_trigger_filtered | irqarray12_trigger[6])) begin
        irqarray12_eventsourceflex198_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex198_clear) begin
            irqarray12_eventsourceflex198_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex198_pending <= irqarray12_eventsourceflex198_pending;
        end
    end
    irqarray12_eventsourceflex199_trigger_d <= irqarray12_interrupts[7];
    if ((irqarray12_eventsourceflex199_trigger_filtered | irqarray12_trigger[7])) begin
        irqarray12_eventsourceflex199_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex199_clear) begin
            irqarray12_eventsourceflex199_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex199_pending <= irqarray12_eventsourceflex199_pending;
        end
    end
    irqarray12_eventsourceflex200_trigger_d <= irqarray12_interrupts[8];
    if ((irqarray12_eventsourceflex200_trigger_filtered | irqarray12_trigger[8])) begin
        irqarray12_eventsourceflex200_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex200_clear) begin
            irqarray12_eventsourceflex200_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex200_pending <= irqarray12_eventsourceflex200_pending;
        end
    end
    irqarray12_eventsourceflex201_trigger_d <= irqarray12_interrupts[9];
    if ((irqarray12_eventsourceflex201_trigger_filtered | irqarray12_trigger[9])) begin
        irqarray12_eventsourceflex201_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex201_clear) begin
            irqarray12_eventsourceflex201_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex201_pending <= irqarray12_eventsourceflex201_pending;
        end
    end
    irqarray12_eventsourceflex202_trigger_d <= irqarray12_interrupts[10];
    if ((irqarray12_eventsourceflex202_trigger_filtered | irqarray12_trigger[10])) begin
        irqarray12_eventsourceflex202_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex202_clear) begin
            irqarray12_eventsourceflex202_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex202_pending <= irqarray12_eventsourceflex202_pending;
        end
    end
    irqarray12_eventsourceflex203_trigger_d <= irqarray12_interrupts[11];
    if ((irqarray12_eventsourceflex203_trigger_filtered | irqarray12_trigger[11])) begin
        irqarray12_eventsourceflex203_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex203_clear) begin
            irqarray12_eventsourceflex203_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex203_pending <= irqarray12_eventsourceflex203_pending;
        end
    end
    irqarray12_eventsourceflex204_trigger_d <= irqarray12_interrupts[12];
    if ((irqarray12_eventsourceflex204_trigger_filtered | irqarray12_trigger[12])) begin
        irqarray12_eventsourceflex204_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex204_clear) begin
            irqarray12_eventsourceflex204_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex204_pending <= irqarray12_eventsourceflex204_pending;
        end
    end
    irqarray12_eventsourceflex205_trigger_d <= irqarray12_interrupts[13];
    if ((irqarray12_eventsourceflex205_trigger_filtered | irqarray12_trigger[13])) begin
        irqarray12_eventsourceflex205_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex205_clear) begin
            irqarray12_eventsourceflex205_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex205_pending <= irqarray12_eventsourceflex205_pending;
        end
    end
    irqarray12_eventsourceflex206_trigger_d <= irqarray12_interrupts[14];
    if ((irqarray12_eventsourceflex206_trigger_filtered | irqarray12_trigger[14])) begin
        irqarray12_eventsourceflex206_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex206_clear) begin
            irqarray12_eventsourceflex206_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex206_pending <= irqarray12_eventsourceflex206_pending;
        end
    end
    irqarray12_eventsourceflex207_trigger_d <= irqarray12_interrupts[15];
    if ((irqarray12_eventsourceflex207_trigger_filtered | irqarray12_trigger[15])) begin
        irqarray12_eventsourceflex207_pending <= 1'd1;
    end else begin
        if (irqarray12_eventsourceflex207_clear) begin
            irqarray12_eventsourceflex207_pending <= 1'd0;
        end else begin
            irqarray12_eventsourceflex207_pending <= irqarray12_eventsourceflex207_pending;
        end
    end
    irqarray13_eventsourceflex208_trigger_d <= irqarray13_interrupts[0];
    if ((irqarray13_eventsourceflex208_trigger_filtered | irqarray13_trigger[0])) begin
        irqarray13_eventsourceflex208_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex208_clear) begin
            irqarray13_eventsourceflex208_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex208_pending <= irqarray13_eventsourceflex208_pending;
        end
    end
    irqarray13_eventsourceflex209_trigger_d <= irqarray13_interrupts[1];
    if ((irqarray13_eventsourceflex209_trigger_filtered | irqarray13_trigger[1])) begin
        irqarray13_eventsourceflex209_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex209_clear) begin
            irqarray13_eventsourceflex209_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex209_pending <= irqarray13_eventsourceflex209_pending;
        end
    end
    irqarray13_eventsourceflex210_trigger_d <= irqarray13_interrupts[2];
    if ((irqarray13_eventsourceflex210_trigger_filtered | irqarray13_trigger[2])) begin
        irqarray13_eventsourceflex210_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex210_clear) begin
            irqarray13_eventsourceflex210_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex210_pending <= irqarray13_eventsourceflex210_pending;
        end
    end
    irqarray13_eventsourceflex211_trigger_d <= irqarray13_interrupts[3];
    if ((irqarray13_eventsourceflex211_trigger_filtered | irqarray13_trigger[3])) begin
        irqarray13_eventsourceflex211_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex211_clear) begin
            irqarray13_eventsourceflex211_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex211_pending <= irqarray13_eventsourceflex211_pending;
        end
    end
    irqarray13_eventsourceflex212_trigger_d <= irqarray13_interrupts[4];
    if ((irqarray13_eventsourceflex212_trigger_filtered | irqarray13_trigger[4])) begin
        irqarray13_eventsourceflex212_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex212_clear) begin
            irqarray13_eventsourceflex212_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex212_pending <= irqarray13_eventsourceflex212_pending;
        end
    end
    irqarray13_eventsourceflex213_trigger_d <= irqarray13_interrupts[5];
    if ((irqarray13_eventsourceflex213_trigger_filtered | irqarray13_trigger[5])) begin
        irqarray13_eventsourceflex213_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex213_clear) begin
            irqarray13_eventsourceflex213_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex213_pending <= irqarray13_eventsourceflex213_pending;
        end
    end
    irqarray13_eventsourceflex214_trigger_d <= irqarray13_interrupts[6];
    if ((irqarray13_eventsourceflex214_trigger_filtered | irqarray13_trigger[6])) begin
        irqarray13_eventsourceflex214_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex214_clear) begin
            irqarray13_eventsourceflex214_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex214_pending <= irqarray13_eventsourceflex214_pending;
        end
    end
    irqarray13_eventsourceflex215_trigger_d <= irqarray13_interrupts[7];
    if ((irqarray13_eventsourceflex215_trigger_filtered | irqarray13_trigger[7])) begin
        irqarray13_eventsourceflex215_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex215_clear) begin
            irqarray13_eventsourceflex215_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex215_pending <= irqarray13_eventsourceflex215_pending;
        end
    end
    irqarray13_eventsourceflex216_trigger_d <= irqarray13_interrupts[8];
    if ((irqarray13_eventsourceflex216_trigger_filtered | irqarray13_trigger[8])) begin
        irqarray13_eventsourceflex216_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex216_clear) begin
            irqarray13_eventsourceflex216_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex216_pending <= irqarray13_eventsourceflex216_pending;
        end
    end
    irqarray13_eventsourceflex217_trigger_d <= irqarray13_interrupts[9];
    if ((irqarray13_eventsourceflex217_trigger_filtered | irqarray13_trigger[9])) begin
        irqarray13_eventsourceflex217_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex217_clear) begin
            irqarray13_eventsourceflex217_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex217_pending <= irqarray13_eventsourceflex217_pending;
        end
    end
    irqarray13_eventsourceflex218_trigger_d <= irqarray13_interrupts[10];
    if ((irqarray13_eventsourceflex218_trigger_filtered | irqarray13_trigger[10])) begin
        irqarray13_eventsourceflex218_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex218_clear) begin
            irqarray13_eventsourceflex218_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex218_pending <= irqarray13_eventsourceflex218_pending;
        end
    end
    irqarray13_eventsourceflex219_trigger_d <= irqarray13_interrupts[11];
    if ((irqarray13_eventsourceflex219_trigger_filtered | irqarray13_trigger[11])) begin
        irqarray13_eventsourceflex219_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex219_clear) begin
            irqarray13_eventsourceflex219_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex219_pending <= irqarray13_eventsourceflex219_pending;
        end
    end
    irqarray13_eventsourceflex220_trigger_d <= irqarray13_interrupts[12];
    if ((irqarray13_eventsourceflex220_trigger_filtered | irqarray13_trigger[12])) begin
        irqarray13_eventsourceflex220_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex220_clear) begin
            irqarray13_eventsourceflex220_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex220_pending <= irqarray13_eventsourceflex220_pending;
        end
    end
    irqarray13_eventsourceflex221_trigger_d <= irqarray13_interrupts[13];
    if ((irqarray13_eventsourceflex221_trigger_filtered | irqarray13_trigger[13])) begin
        irqarray13_eventsourceflex221_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex221_clear) begin
            irqarray13_eventsourceflex221_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex221_pending <= irqarray13_eventsourceflex221_pending;
        end
    end
    irqarray13_eventsourceflex222_trigger_d <= irqarray13_interrupts[14];
    if ((irqarray13_eventsourceflex222_trigger_filtered | irqarray13_trigger[14])) begin
        irqarray13_eventsourceflex222_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex222_clear) begin
            irqarray13_eventsourceflex222_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex222_pending <= irqarray13_eventsourceflex222_pending;
        end
    end
    irqarray13_eventsourceflex223_trigger_d <= irqarray13_interrupts[15];
    if ((irqarray13_eventsourceflex223_trigger_filtered | irqarray13_trigger[15])) begin
        irqarray13_eventsourceflex223_pending <= 1'd1;
    end else begin
        if (irqarray13_eventsourceflex223_clear) begin
            irqarray13_eventsourceflex223_pending <= 1'd0;
        end else begin
            irqarray13_eventsourceflex223_pending <= irqarray13_eventsourceflex223_pending;
        end
    end
    irqarray14_eventsourceflex224_trigger_d <= irqarray14_interrupts[0];
    if ((irqarray14_eventsourceflex224_trigger_filtered | irqarray14_trigger[0])) begin
        irqarray14_eventsourceflex224_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex224_clear) begin
            irqarray14_eventsourceflex224_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex224_pending <= irqarray14_eventsourceflex224_pending;
        end
    end
    irqarray14_eventsourceflex225_trigger_d <= irqarray14_interrupts[1];
    if ((irqarray14_eventsourceflex225_trigger_filtered | irqarray14_trigger[1])) begin
        irqarray14_eventsourceflex225_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex225_clear) begin
            irqarray14_eventsourceflex225_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex225_pending <= irqarray14_eventsourceflex225_pending;
        end
    end
    irqarray14_eventsourceflex226_trigger_d <= irqarray14_interrupts[2];
    if ((irqarray14_eventsourceflex226_trigger_filtered | irqarray14_trigger[2])) begin
        irqarray14_eventsourceflex226_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex226_clear) begin
            irqarray14_eventsourceflex226_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex226_pending <= irqarray14_eventsourceflex226_pending;
        end
    end
    irqarray14_eventsourceflex227_trigger_d <= irqarray14_interrupts[3];
    if ((irqarray14_eventsourceflex227_trigger_filtered | irqarray14_trigger[3])) begin
        irqarray14_eventsourceflex227_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex227_clear) begin
            irqarray14_eventsourceflex227_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex227_pending <= irqarray14_eventsourceflex227_pending;
        end
    end
    irqarray14_eventsourceflex228_trigger_d <= irqarray14_interrupts[4];
    if ((irqarray14_eventsourceflex228_trigger_filtered | irqarray14_trigger[4])) begin
        irqarray14_eventsourceflex228_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex228_clear) begin
            irqarray14_eventsourceflex228_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex228_pending <= irqarray14_eventsourceflex228_pending;
        end
    end
    irqarray14_eventsourceflex229_trigger_d <= irqarray14_interrupts[5];
    if ((irqarray14_eventsourceflex229_trigger_filtered | irqarray14_trigger[5])) begin
        irqarray14_eventsourceflex229_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex229_clear) begin
            irqarray14_eventsourceflex229_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex229_pending <= irqarray14_eventsourceflex229_pending;
        end
    end
    irqarray14_eventsourceflex230_trigger_d <= irqarray14_interrupts[6];
    if ((irqarray14_eventsourceflex230_trigger_filtered | irqarray14_trigger[6])) begin
        irqarray14_eventsourceflex230_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex230_clear) begin
            irqarray14_eventsourceflex230_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex230_pending <= irqarray14_eventsourceflex230_pending;
        end
    end
    irqarray14_eventsourceflex231_trigger_d <= irqarray14_interrupts[7];
    if ((irqarray14_eventsourceflex231_trigger_filtered | irqarray14_trigger[7])) begin
        irqarray14_eventsourceflex231_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex231_clear) begin
            irqarray14_eventsourceflex231_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex231_pending <= irqarray14_eventsourceflex231_pending;
        end
    end
    irqarray14_eventsourceflex232_trigger_d <= irqarray14_interrupts[8];
    if ((irqarray14_eventsourceflex232_trigger_filtered | irqarray14_trigger[8])) begin
        irqarray14_eventsourceflex232_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex232_clear) begin
            irqarray14_eventsourceflex232_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex232_pending <= irqarray14_eventsourceflex232_pending;
        end
    end
    irqarray14_eventsourceflex233_trigger_d <= irqarray14_interrupts[9];
    if ((irqarray14_eventsourceflex233_trigger_filtered | irqarray14_trigger[9])) begin
        irqarray14_eventsourceflex233_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex233_clear) begin
            irqarray14_eventsourceflex233_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex233_pending <= irqarray14_eventsourceflex233_pending;
        end
    end
    irqarray14_eventsourceflex234_trigger_d <= irqarray14_interrupts[10];
    if ((irqarray14_eventsourceflex234_trigger_filtered | irqarray14_trigger[10])) begin
        irqarray14_eventsourceflex234_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex234_clear) begin
            irqarray14_eventsourceflex234_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex234_pending <= irqarray14_eventsourceflex234_pending;
        end
    end
    irqarray14_eventsourceflex235_trigger_d <= irqarray14_interrupts[11];
    if ((irqarray14_eventsourceflex235_trigger_filtered | irqarray14_trigger[11])) begin
        irqarray14_eventsourceflex235_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex235_clear) begin
            irqarray14_eventsourceflex235_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex235_pending <= irqarray14_eventsourceflex235_pending;
        end
    end
    irqarray14_eventsourceflex236_trigger_d <= irqarray14_interrupts[12];
    if ((irqarray14_eventsourceflex236_trigger_filtered | irqarray14_trigger[12])) begin
        irqarray14_eventsourceflex236_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex236_clear) begin
            irqarray14_eventsourceflex236_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex236_pending <= irqarray14_eventsourceflex236_pending;
        end
    end
    irqarray14_eventsourceflex237_trigger_d <= irqarray14_interrupts[13];
    if ((irqarray14_eventsourceflex237_trigger_filtered | irqarray14_trigger[13])) begin
        irqarray14_eventsourceflex237_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex237_clear) begin
            irqarray14_eventsourceflex237_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex237_pending <= irqarray14_eventsourceflex237_pending;
        end
    end
    irqarray14_eventsourceflex238_trigger_d <= irqarray14_interrupts[14];
    if ((irqarray14_eventsourceflex238_trigger_filtered | irqarray14_trigger[14])) begin
        irqarray14_eventsourceflex238_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex238_clear) begin
            irqarray14_eventsourceflex238_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex238_pending <= irqarray14_eventsourceflex238_pending;
        end
    end
    irqarray14_eventsourceflex239_trigger_d <= irqarray14_interrupts[15];
    if ((irqarray14_eventsourceflex239_trigger_filtered | irqarray14_trigger[15])) begin
        irqarray14_eventsourceflex239_pending <= 1'd1;
    end else begin
        if (irqarray14_eventsourceflex239_clear) begin
            irqarray14_eventsourceflex239_pending <= 1'd0;
        end else begin
            irqarray14_eventsourceflex239_pending <= irqarray14_eventsourceflex239_pending;
        end
    end
    irqarray15_eventsourceflex240_trigger_d <= irqarray15_interrupts[0];
    if ((irqarray15_eventsourceflex240_trigger_filtered | irqarray15_trigger[0])) begin
        irqarray15_eventsourceflex240_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex240_clear) begin
            irqarray15_eventsourceflex240_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex240_pending <= irqarray15_eventsourceflex240_pending;
        end
    end
    irqarray15_eventsourceflex241_trigger_d <= irqarray15_interrupts[1];
    if ((irqarray15_eventsourceflex241_trigger_filtered | irqarray15_trigger[1])) begin
        irqarray15_eventsourceflex241_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex241_clear) begin
            irqarray15_eventsourceflex241_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex241_pending <= irqarray15_eventsourceflex241_pending;
        end
    end
    irqarray15_eventsourceflex242_trigger_d <= irqarray15_interrupts[2];
    if ((irqarray15_eventsourceflex242_trigger_filtered | irqarray15_trigger[2])) begin
        irqarray15_eventsourceflex242_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex242_clear) begin
            irqarray15_eventsourceflex242_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex242_pending <= irqarray15_eventsourceflex242_pending;
        end
    end
    irqarray15_eventsourceflex243_trigger_d <= irqarray15_interrupts[3];
    if ((irqarray15_eventsourceflex243_trigger_filtered | irqarray15_trigger[3])) begin
        irqarray15_eventsourceflex243_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex243_clear) begin
            irqarray15_eventsourceflex243_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex243_pending <= irqarray15_eventsourceflex243_pending;
        end
    end
    irqarray15_eventsourceflex244_trigger_d <= irqarray15_interrupts[4];
    if ((irqarray15_eventsourceflex244_trigger_filtered | irqarray15_trigger[4])) begin
        irqarray15_eventsourceflex244_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex244_clear) begin
            irqarray15_eventsourceflex244_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex244_pending <= irqarray15_eventsourceflex244_pending;
        end
    end
    irqarray15_eventsourceflex245_trigger_d <= irqarray15_interrupts[5];
    if ((irqarray15_eventsourceflex245_trigger_filtered | irqarray15_trigger[5])) begin
        irqarray15_eventsourceflex245_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex245_clear) begin
            irqarray15_eventsourceflex245_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex245_pending <= irqarray15_eventsourceflex245_pending;
        end
    end
    irqarray15_eventsourceflex246_trigger_d <= irqarray15_interrupts[6];
    if ((irqarray15_eventsourceflex246_trigger_filtered | irqarray15_trigger[6])) begin
        irqarray15_eventsourceflex246_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex246_clear) begin
            irqarray15_eventsourceflex246_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex246_pending <= irqarray15_eventsourceflex246_pending;
        end
    end
    irqarray15_eventsourceflex247_trigger_d <= irqarray15_interrupts[7];
    if ((irqarray15_eventsourceflex247_trigger_filtered | irqarray15_trigger[7])) begin
        irqarray15_eventsourceflex247_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex247_clear) begin
            irqarray15_eventsourceflex247_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex247_pending <= irqarray15_eventsourceflex247_pending;
        end
    end
    irqarray15_eventsourceflex248_trigger_d <= irqarray15_interrupts[8];
    if ((irqarray15_eventsourceflex248_trigger_filtered | irqarray15_trigger[8])) begin
        irqarray15_eventsourceflex248_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex248_clear) begin
            irqarray15_eventsourceflex248_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex248_pending <= irqarray15_eventsourceflex248_pending;
        end
    end
    irqarray15_eventsourceflex249_trigger_d <= irqarray15_interrupts[9];
    if ((irqarray15_eventsourceflex249_trigger_filtered | irqarray15_trigger[9])) begin
        irqarray15_eventsourceflex249_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex249_clear) begin
            irqarray15_eventsourceflex249_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex249_pending <= irqarray15_eventsourceflex249_pending;
        end
    end
    irqarray15_eventsourceflex250_trigger_d <= irqarray15_interrupts[10];
    if ((irqarray15_eventsourceflex250_trigger_filtered | irqarray15_trigger[10])) begin
        irqarray15_eventsourceflex250_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex250_clear) begin
            irqarray15_eventsourceflex250_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex250_pending <= irqarray15_eventsourceflex250_pending;
        end
    end
    irqarray15_eventsourceflex251_trigger_d <= irqarray15_interrupts[11];
    if ((irqarray15_eventsourceflex251_trigger_filtered | irqarray15_trigger[11])) begin
        irqarray15_eventsourceflex251_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex251_clear) begin
            irqarray15_eventsourceflex251_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex251_pending <= irqarray15_eventsourceflex251_pending;
        end
    end
    irqarray15_eventsourceflex252_trigger_d <= irqarray15_interrupts[12];
    if ((irqarray15_eventsourceflex252_trigger_filtered | irqarray15_trigger[12])) begin
        irqarray15_eventsourceflex252_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex252_clear) begin
            irqarray15_eventsourceflex252_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex252_pending <= irqarray15_eventsourceflex252_pending;
        end
    end
    irqarray15_eventsourceflex253_trigger_d <= irqarray15_interrupts[13];
    if ((irqarray15_eventsourceflex253_trigger_filtered | irqarray15_trigger[13])) begin
        irqarray15_eventsourceflex253_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex253_clear) begin
            irqarray15_eventsourceflex253_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex253_pending <= irqarray15_eventsourceflex253_pending;
        end
    end
    irqarray15_eventsourceflex254_trigger_d <= irqarray15_interrupts[14];
    if ((irqarray15_eventsourceflex254_trigger_filtered | irqarray15_trigger[14])) begin
        irqarray15_eventsourceflex254_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex254_clear) begin
            irqarray15_eventsourceflex254_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex254_pending <= irqarray15_eventsourceflex254_pending;
        end
    end
    irqarray15_eventsourceflex255_trigger_d <= irqarray15_interrupts[15];
    if ((irqarray15_eventsourceflex255_trigger_filtered | irqarray15_trigger[15])) begin
        irqarray15_eventsourceflex255_pending <= 1'd1;
    end else begin
        if (irqarray15_eventsourceflex255_clear) begin
            irqarray15_eventsourceflex255_pending <= 1'd0;
        end else begin
            irqarray15_eventsourceflex255_pending <= irqarray15_eventsourceflex255_pending;
        end
    end
    irqarray16_eventsourceflex256_trigger_d <= irqarray16_interrupts[0];
    if ((irqarray16_eventsourceflex256_trigger_filtered | irqarray16_trigger[0])) begin
        irqarray16_eventsourceflex256_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex256_clear) begin
            irqarray16_eventsourceflex256_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex256_pending <= irqarray16_eventsourceflex256_pending;
        end
    end
    irqarray16_eventsourceflex257_trigger_d <= irqarray16_interrupts[1];
    if ((irqarray16_eventsourceflex257_trigger_filtered | irqarray16_trigger[1])) begin
        irqarray16_eventsourceflex257_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex257_clear) begin
            irqarray16_eventsourceflex257_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex257_pending <= irqarray16_eventsourceflex257_pending;
        end
    end
    irqarray16_eventsourceflex258_trigger_d <= irqarray16_interrupts[2];
    if ((irqarray16_eventsourceflex258_trigger_filtered | irqarray16_trigger[2])) begin
        irqarray16_eventsourceflex258_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex258_clear) begin
            irqarray16_eventsourceflex258_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex258_pending <= irqarray16_eventsourceflex258_pending;
        end
    end
    irqarray16_eventsourceflex259_trigger_d <= irqarray16_interrupts[3];
    if ((irqarray16_eventsourceflex259_trigger_filtered | irqarray16_trigger[3])) begin
        irqarray16_eventsourceflex259_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex259_clear) begin
            irqarray16_eventsourceflex259_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex259_pending <= irqarray16_eventsourceflex259_pending;
        end
    end
    irqarray16_eventsourceflex260_trigger_d <= irqarray16_interrupts[4];
    if ((irqarray16_eventsourceflex260_trigger_filtered | irqarray16_trigger[4])) begin
        irqarray16_eventsourceflex260_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex260_clear) begin
            irqarray16_eventsourceflex260_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex260_pending <= irqarray16_eventsourceflex260_pending;
        end
    end
    irqarray16_eventsourceflex261_trigger_d <= irqarray16_interrupts[5];
    if ((irqarray16_eventsourceflex261_trigger_filtered | irqarray16_trigger[5])) begin
        irqarray16_eventsourceflex261_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex261_clear) begin
            irqarray16_eventsourceflex261_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex261_pending <= irqarray16_eventsourceflex261_pending;
        end
    end
    irqarray16_eventsourceflex262_trigger_d <= irqarray16_interrupts[6];
    if ((irqarray16_eventsourceflex262_trigger_filtered | irqarray16_trigger[6])) begin
        irqarray16_eventsourceflex262_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex262_clear) begin
            irqarray16_eventsourceflex262_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex262_pending <= irqarray16_eventsourceflex262_pending;
        end
    end
    irqarray16_eventsourceflex263_trigger_d <= irqarray16_interrupts[7];
    if ((irqarray16_eventsourceflex263_trigger_filtered | irqarray16_trigger[7])) begin
        irqarray16_eventsourceflex263_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex263_clear) begin
            irqarray16_eventsourceflex263_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex263_pending <= irqarray16_eventsourceflex263_pending;
        end
    end
    irqarray16_eventsourceflex264_trigger_d <= irqarray16_interrupts[8];
    if ((irqarray16_eventsourceflex264_trigger_filtered | irqarray16_trigger[8])) begin
        irqarray16_eventsourceflex264_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex264_clear) begin
            irqarray16_eventsourceflex264_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex264_pending <= irqarray16_eventsourceflex264_pending;
        end
    end
    irqarray16_eventsourceflex265_trigger_d <= irqarray16_interrupts[9];
    if ((irqarray16_eventsourceflex265_trigger_filtered | irqarray16_trigger[9])) begin
        irqarray16_eventsourceflex265_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex265_clear) begin
            irqarray16_eventsourceflex265_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex265_pending <= irqarray16_eventsourceflex265_pending;
        end
    end
    irqarray16_eventsourceflex266_trigger_d <= irqarray16_interrupts[10];
    if ((irqarray16_eventsourceflex266_trigger_filtered | irqarray16_trigger[10])) begin
        irqarray16_eventsourceflex266_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex266_clear) begin
            irqarray16_eventsourceflex266_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex266_pending <= irqarray16_eventsourceflex266_pending;
        end
    end
    irqarray16_eventsourceflex267_trigger_d <= irqarray16_interrupts[11];
    if ((irqarray16_eventsourceflex267_trigger_filtered | irqarray16_trigger[11])) begin
        irqarray16_eventsourceflex267_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex267_clear) begin
            irqarray16_eventsourceflex267_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex267_pending <= irqarray16_eventsourceflex267_pending;
        end
    end
    irqarray16_eventsourceflex268_trigger_d <= irqarray16_interrupts[12];
    if ((irqarray16_eventsourceflex268_trigger_filtered | irqarray16_trigger[12])) begin
        irqarray16_eventsourceflex268_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex268_clear) begin
            irqarray16_eventsourceflex268_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex268_pending <= irqarray16_eventsourceflex268_pending;
        end
    end
    irqarray16_eventsourceflex269_trigger_d <= irqarray16_interrupts[13];
    if ((irqarray16_eventsourceflex269_trigger_filtered | irqarray16_trigger[13])) begin
        irqarray16_eventsourceflex269_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex269_clear) begin
            irqarray16_eventsourceflex269_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex269_pending <= irqarray16_eventsourceflex269_pending;
        end
    end
    irqarray16_eventsourceflex270_trigger_d <= irqarray16_interrupts[14];
    if ((irqarray16_eventsourceflex270_trigger_filtered | irqarray16_trigger[14])) begin
        irqarray16_eventsourceflex270_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex270_clear) begin
            irqarray16_eventsourceflex270_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex270_pending <= irqarray16_eventsourceflex270_pending;
        end
    end
    irqarray16_eventsourceflex271_trigger_d <= irqarray16_interrupts[15];
    if ((irqarray16_eventsourceflex271_trigger_filtered | irqarray16_trigger[15])) begin
        irqarray16_eventsourceflex271_pending <= 1'd1;
    end else begin
        if (irqarray16_eventsourceflex271_clear) begin
            irqarray16_eventsourceflex271_pending <= 1'd0;
        end else begin
            irqarray16_eventsourceflex271_pending <= irqarray16_eventsourceflex271_pending;
        end
    end
    irqarray17_eventsourceflex272_trigger_d <= irqarray17_interrupts[0];
    if ((irqarray17_eventsourceflex272_trigger_filtered | irqarray17_trigger[0])) begin
        irqarray17_eventsourceflex272_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex272_clear) begin
            irqarray17_eventsourceflex272_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex272_pending <= irqarray17_eventsourceflex272_pending;
        end
    end
    irqarray17_eventsourceflex273_trigger_d <= irqarray17_interrupts[1];
    if ((irqarray17_eventsourceflex273_trigger_filtered | irqarray17_trigger[1])) begin
        irqarray17_eventsourceflex273_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex273_clear) begin
            irqarray17_eventsourceflex273_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex273_pending <= irqarray17_eventsourceflex273_pending;
        end
    end
    irqarray17_eventsourceflex274_trigger_d <= irqarray17_interrupts[2];
    if ((irqarray17_eventsourceflex274_trigger_filtered | irqarray17_trigger[2])) begin
        irqarray17_eventsourceflex274_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex274_clear) begin
            irqarray17_eventsourceflex274_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex274_pending <= irqarray17_eventsourceflex274_pending;
        end
    end
    irqarray17_eventsourceflex275_trigger_d <= irqarray17_interrupts[3];
    if ((irqarray17_eventsourceflex275_trigger_filtered | irqarray17_trigger[3])) begin
        irqarray17_eventsourceflex275_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex275_clear) begin
            irqarray17_eventsourceflex275_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex275_pending <= irqarray17_eventsourceflex275_pending;
        end
    end
    irqarray17_eventsourceflex276_trigger_d <= irqarray17_interrupts[4];
    if ((irqarray17_eventsourceflex276_trigger_filtered | irqarray17_trigger[4])) begin
        irqarray17_eventsourceflex276_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex276_clear) begin
            irqarray17_eventsourceflex276_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex276_pending <= irqarray17_eventsourceflex276_pending;
        end
    end
    irqarray17_eventsourceflex277_trigger_d <= irqarray17_interrupts[5];
    if ((irqarray17_eventsourceflex277_trigger_filtered | irqarray17_trigger[5])) begin
        irqarray17_eventsourceflex277_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex277_clear) begin
            irqarray17_eventsourceflex277_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex277_pending <= irqarray17_eventsourceflex277_pending;
        end
    end
    irqarray17_eventsourceflex278_trigger_d <= irqarray17_interrupts[6];
    if ((irqarray17_eventsourceflex278_trigger_filtered | irqarray17_trigger[6])) begin
        irqarray17_eventsourceflex278_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex278_clear) begin
            irqarray17_eventsourceflex278_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex278_pending <= irqarray17_eventsourceflex278_pending;
        end
    end
    irqarray17_eventsourceflex279_trigger_d <= irqarray17_interrupts[7];
    if ((irqarray17_eventsourceflex279_trigger_filtered | irqarray17_trigger[7])) begin
        irqarray17_eventsourceflex279_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex279_clear) begin
            irqarray17_eventsourceflex279_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex279_pending <= irqarray17_eventsourceflex279_pending;
        end
    end
    irqarray17_eventsourceflex280_trigger_d <= irqarray17_interrupts[8];
    if ((irqarray17_eventsourceflex280_trigger_filtered | irqarray17_trigger[8])) begin
        irqarray17_eventsourceflex280_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex280_clear) begin
            irqarray17_eventsourceflex280_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex280_pending <= irqarray17_eventsourceflex280_pending;
        end
    end
    irqarray17_eventsourceflex281_trigger_d <= irqarray17_interrupts[9];
    if ((irqarray17_eventsourceflex281_trigger_filtered | irqarray17_trigger[9])) begin
        irqarray17_eventsourceflex281_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex281_clear) begin
            irqarray17_eventsourceflex281_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex281_pending <= irqarray17_eventsourceflex281_pending;
        end
    end
    irqarray17_eventsourceflex282_trigger_d <= irqarray17_interrupts[10];
    if ((irqarray17_eventsourceflex282_trigger_filtered | irqarray17_trigger[10])) begin
        irqarray17_eventsourceflex282_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex282_clear) begin
            irqarray17_eventsourceflex282_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex282_pending <= irqarray17_eventsourceflex282_pending;
        end
    end
    irqarray17_eventsourceflex283_trigger_d <= irqarray17_interrupts[11];
    if ((irqarray17_eventsourceflex283_trigger_filtered | irqarray17_trigger[11])) begin
        irqarray17_eventsourceflex283_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex283_clear) begin
            irqarray17_eventsourceflex283_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex283_pending <= irqarray17_eventsourceflex283_pending;
        end
    end
    irqarray17_eventsourceflex284_trigger_d <= irqarray17_interrupts[12];
    if ((irqarray17_eventsourceflex284_trigger_filtered | irqarray17_trigger[12])) begin
        irqarray17_eventsourceflex284_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex284_clear) begin
            irqarray17_eventsourceflex284_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex284_pending <= irqarray17_eventsourceflex284_pending;
        end
    end
    irqarray17_eventsourceflex285_trigger_d <= irqarray17_interrupts[13];
    if ((irqarray17_eventsourceflex285_trigger_filtered | irqarray17_trigger[13])) begin
        irqarray17_eventsourceflex285_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex285_clear) begin
            irqarray17_eventsourceflex285_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex285_pending <= irqarray17_eventsourceflex285_pending;
        end
    end
    irqarray17_eventsourceflex286_trigger_d <= irqarray17_interrupts[14];
    if ((irqarray17_eventsourceflex286_trigger_filtered | irqarray17_trigger[14])) begin
        irqarray17_eventsourceflex286_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex286_clear) begin
            irqarray17_eventsourceflex286_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex286_pending <= irqarray17_eventsourceflex286_pending;
        end
    end
    irqarray17_eventsourceflex287_trigger_d <= irqarray17_interrupts[15];
    if ((irqarray17_eventsourceflex287_trigger_filtered | irqarray17_trigger[15])) begin
        irqarray17_eventsourceflex287_pending <= 1'd1;
    end else begin
        if (irqarray17_eventsourceflex287_clear) begin
            irqarray17_eventsourceflex287_pending <= 1'd0;
        end else begin
            irqarray17_eventsourceflex287_pending <= irqarray17_eventsourceflex287_pending;
        end
    end
    irqarray18_eventsourceflex288_trigger_d <= irqarray18_interrupts[0];
    if ((irqarray18_eventsourceflex288_trigger_filtered | irqarray18_trigger[0])) begin
        irqarray18_eventsourceflex288_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex288_clear) begin
            irqarray18_eventsourceflex288_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex288_pending <= irqarray18_eventsourceflex288_pending;
        end
    end
    irqarray18_eventsourceflex289_trigger_d <= irqarray18_interrupts[1];
    if ((irqarray18_eventsourceflex289_trigger_filtered | irqarray18_trigger[1])) begin
        irqarray18_eventsourceflex289_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex289_clear) begin
            irqarray18_eventsourceflex289_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex289_pending <= irqarray18_eventsourceflex289_pending;
        end
    end
    irqarray18_eventsourceflex290_trigger_d <= irqarray18_interrupts[2];
    if ((irqarray18_eventsourceflex290_trigger_filtered | irqarray18_trigger[2])) begin
        irqarray18_eventsourceflex290_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex290_clear) begin
            irqarray18_eventsourceflex290_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex290_pending <= irqarray18_eventsourceflex290_pending;
        end
    end
    irqarray18_eventsourceflex291_trigger_d <= irqarray18_interrupts[3];
    if ((irqarray18_eventsourceflex291_trigger_filtered | irqarray18_trigger[3])) begin
        irqarray18_eventsourceflex291_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex291_clear) begin
            irqarray18_eventsourceflex291_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex291_pending <= irqarray18_eventsourceflex291_pending;
        end
    end
    irqarray18_eventsourceflex292_trigger_d <= irqarray18_interrupts[4];
    if ((irqarray18_eventsourceflex292_trigger_filtered | irqarray18_trigger[4])) begin
        irqarray18_eventsourceflex292_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex292_clear) begin
            irqarray18_eventsourceflex292_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex292_pending <= irqarray18_eventsourceflex292_pending;
        end
    end
    irqarray18_eventsourceflex293_trigger_d <= irqarray18_interrupts[5];
    if ((irqarray18_eventsourceflex293_trigger_filtered | irqarray18_trigger[5])) begin
        irqarray18_eventsourceflex293_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex293_clear) begin
            irqarray18_eventsourceflex293_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex293_pending <= irqarray18_eventsourceflex293_pending;
        end
    end
    irqarray18_eventsourceflex294_trigger_d <= irqarray18_interrupts[6];
    if ((irqarray18_eventsourceflex294_trigger_filtered | irqarray18_trigger[6])) begin
        irqarray18_eventsourceflex294_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex294_clear) begin
            irqarray18_eventsourceflex294_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex294_pending <= irqarray18_eventsourceflex294_pending;
        end
    end
    irqarray18_eventsourceflex295_trigger_d <= irqarray18_interrupts[7];
    if ((irqarray18_eventsourceflex295_trigger_filtered | irqarray18_trigger[7])) begin
        irqarray18_eventsourceflex295_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex295_clear) begin
            irqarray18_eventsourceflex295_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex295_pending <= irqarray18_eventsourceflex295_pending;
        end
    end
    irqarray18_eventsourceflex296_trigger_d <= irqarray18_interrupts[8];
    if ((irqarray18_eventsourceflex296_trigger_filtered | irqarray18_trigger[8])) begin
        irqarray18_eventsourceflex296_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex296_clear) begin
            irqarray18_eventsourceflex296_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex296_pending <= irqarray18_eventsourceflex296_pending;
        end
    end
    irqarray18_eventsourceflex297_trigger_d <= irqarray18_interrupts[9];
    if ((irqarray18_eventsourceflex297_trigger_filtered | irqarray18_trigger[9])) begin
        irqarray18_eventsourceflex297_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex297_clear) begin
            irqarray18_eventsourceflex297_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex297_pending <= irqarray18_eventsourceflex297_pending;
        end
    end
    irqarray18_eventsourceflex298_trigger_d <= irqarray18_interrupts[10];
    if ((irqarray18_eventsourceflex298_trigger_filtered | irqarray18_trigger[10])) begin
        irqarray18_eventsourceflex298_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex298_clear) begin
            irqarray18_eventsourceflex298_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex298_pending <= irqarray18_eventsourceflex298_pending;
        end
    end
    irqarray18_eventsourceflex299_trigger_d <= irqarray18_interrupts[11];
    if ((irqarray18_eventsourceflex299_trigger_filtered | irqarray18_trigger[11])) begin
        irqarray18_eventsourceflex299_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex299_clear) begin
            irqarray18_eventsourceflex299_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex299_pending <= irqarray18_eventsourceflex299_pending;
        end
    end
    irqarray18_eventsourceflex300_trigger_d <= irqarray18_interrupts[12];
    if ((irqarray18_eventsourceflex300_trigger_filtered | irqarray18_trigger[12])) begin
        irqarray18_eventsourceflex300_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex300_clear) begin
            irqarray18_eventsourceflex300_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex300_pending <= irqarray18_eventsourceflex300_pending;
        end
    end
    irqarray18_eventsourceflex301_trigger_d <= irqarray18_interrupts[13];
    if ((irqarray18_eventsourceflex301_trigger_filtered | irqarray18_trigger[13])) begin
        irqarray18_eventsourceflex301_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex301_clear) begin
            irqarray18_eventsourceflex301_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex301_pending <= irqarray18_eventsourceflex301_pending;
        end
    end
    irqarray18_eventsourceflex302_trigger_d <= irqarray18_interrupts[14];
    if ((irqarray18_eventsourceflex302_trigger_filtered | irqarray18_trigger[14])) begin
        irqarray18_eventsourceflex302_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex302_clear) begin
            irqarray18_eventsourceflex302_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex302_pending <= irqarray18_eventsourceflex302_pending;
        end
    end
    irqarray18_eventsourceflex303_trigger_d <= irqarray18_interrupts[15];
    if ((irqarray18_eventsourceflex303_trigger_filtered | irqarray18_trigger[15])) begin
        irqarray18_eventsourceflex303_pending <= 1'd1;
    end else begin
        if (irqarray18_eventsourceflex303_clear) begin
            irqarray18_eventsourceflex303_pending <= 1'd0;
        end else begin
            irqarray18_eventsourceflex303_pending <= irqarray18_eventsourceflex303_pending;
        end
    end
    irqarray19_eventsourceflex304_trigger_d <= irqarray19_interrupts[0];
    if ((irqarray19_eventsourceflex304_trigger_filtered | irqarray19_trigger[0])) begin
        irqarray19_eventsourceflex304_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex304_clear) begin
            irqarray19_eventsourceflex304_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex304_pending <= irqarray19_eventsourceflex304_pending;
        end
    end
    irqarray19_eventsourceflex305_trigger_d <= irqarray19_interrupts[1];
    if ((irqarray19_eventsourceflex305_trigger_filtered | irqarray19_trigger[1])) begin
        irqarray19_eventsourceflex305_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex305_clear) begin
            irqarray19_eventsourceflex305_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex305_pending <= irqarray19_eventsourceflex305_pending;
        end
    end
    irqarray19_eventsourceflex306_trigger_d <= irqarray19_interrupts[2];
    if ((irqarray19_eventsourceflex306_trigger_filtered | irqarray19_trigger[2])) begin
        irqarray19_eventsourceflex306_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex306_clear) begin
            irqarray19_eventsourceflex306_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex306_pending <= irqarray19_eventsourceflex306_pending;
        end
    end
    irqarray19_eventsourceflex307_trigger_d <= irqarray19_interrupts[3];
    if ((irqarray19_eventsourceflex307_trigger_filtered | irqarray19_trigger[3])) begin
        irqarray19_eventsourceflex307_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex307_clear) begin
            irqarray19_eventsourceflex307_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex307_pending <= irqarray19_eventsourceflex307_pending;
        end
    end
    irqarray19_eventsourceflex308_trigger_d <= irqarray19_interrupts[4];
    if ((irqarray19_eventsourceflex308_trigger_filtered | irqarray19_trigger[4])) begin
        irqarray19_eventsourceflex308_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex308_clear) begin
            irqarray19_eventsourceflex308_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex308_pending <= irqarray19_eventsourceflex308_pending;
        end
    end
    irqarray19_eventsourceflex309_trigger_d <= irqarray19_interrupts[5];
    if ((irqarray19_eventsourceflex309_trigger_filtered | irqarray19_trigger[5])) begin
        irqarray19_eventsourceflex309_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex309_clear) begin
            irqarray19_eventsourceflex309_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex309_pending <= irqarray19_eventsourceflex309_pending;
        end
    end
    irqarray19_eventsourceflex310_trigger_d <= irqarray19_interrupts[6];
    if ((irqarray19_eventsourceflex310_trigger_filtered | irqarray19_trigger[6])) begin
        irqarray19_eventsourceflex310_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex310_clear) begin
            irqarray19_eventsourceflex310_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex310_pending <= irqarray19_eventsourceflex310_pending;
        end
    end
    irqarray19_eventsourceflex311_trigger_d <= irqarray19_interrupts[7];
    if ((irqarray19_eventsourceflex311_trigger_filtered | irqarray19_trigger[7])) begin
        irqarray19_eventsourceflex311_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex311_clear) begin
            irqarray19_eventsourceflex311_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex311_pending <= irqarray19_eventsourceflex311_pending;
        end
    end
    irqarray19_eventsourceflex312_trigger_d <= irqarray19_interrupts[8];
    if ((irqarray19_eventsourceflex312_trigger_filtered | irqarray19_trigger[8])) begin
        irqarray19_eventsourceflex312_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex312_clear) begin
            irqarray19_eventsourceflex312_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex312_pending <= irqarray19_eventsourceflex312_pending;
        end
    end
    irqarray19_eventsourceflex313_trigger_d <= irqarray19_interrupts[9];
    if ((irqarray19_eventsourceflex313_trigger_filtered | irqarray19_trigger[9])) begin
        irqarray19_eventsourceflex313_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex313_clear) begin
            irqarray19_eventsourceflex313_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex313_pending <= irqarray19_eventsourceflex313_pending;
        end
    end
    irqarray19_eventsourceflex314_trigger_d <= irqarray19_interrupts[10];
    if ((irqarray19_eventsourceflex314_trigger_filtered | irqarray19_trigger[10])) begin
        irqarray19_eventsourceflex314_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex314_clear) begin
            irqarray19_eventsourceflex314_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex314_pending <= irqarray19_eventsourceflex314_pending;
        end
    end
    irqarray19_eventsourceflex315_trigger_d <= irqarray19_interrupts[11];
    if ((irqarray19_eventsourceflex315_trigger_filtered | irqarray19_trigger[11])) begin
        irqarray19_eventsourceflex315_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex315_clear) begin
            irqarray19_eventsourceflex315_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex315_pending <= irqarray19_eventsourceflex315_pending;
        end
    end
    irqarray19_eventsourceflex316_trigger_d <= irqarray19_interrupts[12];
    if ((irqarray19_eventsourceflex316_trigger_filtered | irqarray19_trigger[12])) begin
        irqarray19_eventsourceflex316_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex316_clear) begin
            irqarray19_eventsourceflex316_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex316_pending <= irqarray19_eventsourceflex316_pending;
        end
    end
    irqarray19_eventsourceflex317_trigger_d <= irqarray19_interrupts[13];
    if ((irqarray19_eventsourceflex317_trigger_filtered | irqarray19_trigger[13])) begin
        irqarray19_eventsourceflex317_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex317_clear) begin
            irqarray19_eventsourceflex317_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex317_pending <= irqarray19_eventsourceflex317_pending;
        end
    end
    irqarray19_eventsourceflex318_trigger_d <= irqarray19_interrupts[14];
    if ((irqarray19_eventsourceflex318_trigger_filtered | irqarray19_trigger[14])) begin
        irqarray19_eventsourceflex318_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex318_clear) begin
            irqarray19_eventsourceflex318_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex318_pending <= irqarray19_eventsourceflex318_pending;
        end
    end
    irqarray19_eventsourceflex319_trigger_d <= irqarray19_interrupts[15];
    if ((irqarray19_eventsourceflex319_trigger_filtered | irqarray19_trigger[15])) begin
        irqarray19_eventsourceflex319_pending <= 1'd1;
    end else begin
        if (irqarray19_eventsourceflex319_clear) begin
            irqarray19_eventsourceflex319_pending <= 1'd0;
        end else begin
            irqarray19_eventsourceflex319_pending <= irqarray19_eventsourceflex319_pending;
        end
    end
    if (ticktimer_reset_xfer_o) begin
        ticktimer_timer0 <= 1'd0;
        ticktimer_prescaler <= ticktimer_clkspertick;
    end else begin
        if (ticktimer_load_xfer_o) begin
            ticktimer_prescaler <= ticktimer_clkspertick;
            ticktimer_timer0 <= ticktimer_resume_sync_o;
        end else begin
            if ((ticktimer_prescaler == 1'd0)) begin
                ticktimer_prescaler <= ticktimer_clkspertick;
                if ((ticktimer_pause1 == 1'd0)) begin
                    ticktimer_timer0 <= (ticktimer_timer0 + 1'd1);
                    ticktimer_paused1 <= 1'd0;
                end else begin
                    ticktimer_timer0 <= ticktimer_timer0;
                    ticktimer_paused1 <= 1'd1;
                end
            end else begin
                ticktimer_prescaler <= (ticktimer_prescaler - 1'd1);
            end
        end
    end
    ticktimer_alarm3 <= (ticktimer_target_xfer_o <= ticktimer_timer0);
    ticktimer_load_xfer_ps_toggle_o_r <= ticktimer_load_xfer_ps_toggle_o;
    if (ticktimer_load_xfer_ps_ack_i) begin
        ticktimer_load_xfer_ps_ack_toggle_i <= (~ticktimer_load_xfer_ps_ack_toggle_i);
    end
    ticktimer_timer_sync_starter <= 1'd0;
    if (ticktimer_timer_sync_pong_o) begin
        ticktimer_timer_sync_ibuffer <= ticktimer_timer_sync_i;
    end
    if (ticktimer_timer_sync_ping_i) begin
        ticktimer_timer_sync_ping_toggle_i <= (~ticktimer_timer_sync_ping_toggle_i);
    end
    ticktimer_timer_sync_pong_toggle_o_r <= ticktimer_timer_sync_pong_toggle_o;
    if (ticktimer_timer_sync_wait) begin
        if ((~ticktimer_timer_sync_done)) begin
            ticktimer_timer_sync_count <= (ticktimer_timer_sync_count - 1'd1);
        end
    end else begin
        ticktimer_timer_sync_count <= 8'd128;
    end
    ticktimer_resume_sync_ping_o1 <= ticktimer_resume_sync_ping_o0;
    if (ticktimer_resume_sync_ping_o1) begin
        ticktimer_resume_sync_o <= ticktimer_resume_sync_obuffer;
    end
    ticktimer_resume_sync_ping_toggle_o_r <= ticktimer_resume_sync_ping_toggle_o;
    if (ticktimer_resume_sync_pong_i) begin
        ticktimer_resume_sync_pong_toggle_i <= (~ticktimer_resume_sync_pong_toggle_i);
    end
    ticktimer_reset_xfer_ps_toggle_o_r <= ticktimer_reset_xfer_ps_toggle_o;
    if (ticktimer_reset_xfer_ps_ack_i) begin
        ticktimer_reset_xfer_ps_ack_toggle_i <= (~ticktimer_reset_xfer_ps_ack_toggle_i);
    end
    ticktimer_ping_ps_toggle_o_r <= ticktimer_ping_ps_toggle_o;
    if (ticktimer_ping_ps_ack_i) begin
        ticktimer_ping_ps_ack_toggle_i <= (~ticktimer_ping_ps_ack_toggle_i);
    end
    if (ticktimer_pong_i) begin
        ticktimer_pong_blind <= 1'd1;
    end
    if (ticktimer_pong_ps_ack_o) begin
        ticktimer_pong_blind <= 1'd0;
    end
    if (ticktimer_pong_ps_i) begin
        ticktimer_pong_ps_toggle_i <= (~ticktimer_pong_ps_toggle_i);
    end
    ticktimer_pong_ps_ack_toggle_o_r <= ticktimer_pong_ps_ack_toggle_o;
    ticktimer_target_xfer_ping_o1 <= ticktimer_target_xfer_ping_o0;
    if (ticktimer_target_xfer_ping_o1) begin
        ticktimer_target_xfer_o <= ticktimer_target_xfer_obuffer;
    end
    ticktimer_target_xfer_ping_toggle_o_r <= ticktimer_target_xfer_ping_toggle_o;
    if (ticktimer_target_xfer_pong_i) begin
        ticktimer_target_xfer_pong_toggle_i <= (~ticktimer_target_xfer_pong_toggle_i);
    end
    if (ticktimer_msleep_target_re) begin
        ticktimer_lockout_alarm <= 1'd1;
    end else begin
        if (ticktimer_pong_o) begin
            ticktimer_lockout_alarm <= 1'd0;
        end else begin
            ticktimer_lockout_alarm <= ticktimer_lockout_alarm;
        end
    end
    if (ticktimer_load_xfer_i) begin
        ticktimer_load_xfer_blind <= 1'd1;
    end
    if (ticktimer_load_xfer_ps_ack_o) begin
        ticktimer_load_xfer_blind <= 1'd0;
    end
    if (ticktimer_load_xfer_ps_i) begin
        ticktimer_load_xfer_ps_toggle_i <= (~ticktimer_load_xfer_ps_toggle_i);
    end
    ticktimer_load_xfer_ps_ack_toggle_o_r <= ticktimer_load_xfer_ps_ack_toggle_o;
    ticktimer_timer_sync_ping_o1 <= ticktimer_timer_sync_ping_o0;
    if (ticktimer_timer_sync_ping_o1) begin
        ticktimer_timer_sync_o <= ticktimer_timer_sync_obuffer;
    end
    ticktimer_timer_sync_ping_toggle_o_r <= ticktimer_timer_sync_ping_toggle_o;
    if (ticktimer_timer_sync_pong_i) begin
        ticktimer_timer_sync_pong_toggle_i <= (~ticktimer_timer_sync_pong_toggle_i);
    end
    ticktimer_resume_sync_starter <= 1'd0;
    if (ticktimer_resume_sync_pong_o) begin
        ticktimer_resume_sync_ibuffer <= ticktimer_resume_sync_i;
    end
    if (ticktimer_resume_sync_ping_i) begin
        ticktimer_resume_sync_ping_toggle_i <= (~ticktimer_resume_sync_ping_toggle_i);
    end
    ticktimer_resume_sync_pong_toggle_o_r <= ticktimer_resume_sync_pong_toggle_o;
    if (ticktimer_resume_sync_wait) begin
        if ((~ticktimer_resume_sync_done)) begin
            ticktimer_resume_sync_count <= (ticktimer_resume_sync_count - 1'd1);
        end
    end else begin
        ticktimer_resume_sync_count <= 8'd128;
    end
    if (ticktimer_reset_xfer_i) begin
        ticktimer_reset_xfer_blind <= 1'd1;
    end
    if (ticktimer_reset_xfer_ps_ack_o) begin
        ticktimer_reset_xfer_blind <= 1'd0;
    end
    if (ticktimer_reset_xfer_ps_i) begin
        ticktimer_reset_xfer_ps_toggle_i <= (~ticktimer_reset_xfer_ps_toggle_i);
    end
    ticktimer_reset_xfer_ps_ack_toggle_o_r <= ticktimer_reset_xfer_ps_ack_toggle_o;
    if (ticktimer_ping_i) begin
        ticktimer_ping_blind <= 1'd1;
    end
    if (ticktimer_ping_ps_ack_o) begin
        ticktimer_ping_blind <= 1'd0;
    end
    if (ticktimer_ping_ps_i) begin
        ticktimer_ping_ps_toggle_i <= (~ticktimer_ping_ps_toggle_i);
    end
    ticktimer_ping_ps_ack_toggle_o_r <= ticktimer_ping_ps_ack_toggle_o;
    ticktimer_pong_ps_toggle_o_r <= ticktimer_pong_ps_toggle_o;
    if (ticktimer_pong_ps_ack_i) begin
        ticktimer_pong_ps_ack_toggle_i <= (~ticktimer_pong_ps_ack_toggle_i);
    end
    ticktimer_target_xfer_starter <= 1'd0;
    if (ticktimer_target_xfer_pong_o) begin
        ticktimer_target_xfer_ibuffer <= ticktimer_target_xfer_i;
    end
    if (ticktimer_target_xfer_ping_i) begin
        ticktimer_target_xfer_ping_toggle_i <= (~ticktimer_target_xfer_ping_toggle_i);
    end
    ticktimer_target_xfer_pong_toggle_o_r <= ticktimer_target_xfer_pong_toggle_o;
    if (ticktimer_target_xfer_wait) begin
        if ((~ticktimer_target_xfer_done)) begin
            ticktimer_target_xfer_count <= (ticktimer_target_xfer_count - 1'd1);
        end
    end else begin
        ticktimer_target_xfer_count <= 8'd128;
    end
    if ((d11ctime_counter == 1'd0)) begin
        d11ctime_counter <= d11ctime_count;
        d11ctime_heartbeat <= (~d11ctime_heartbeat);
    end else begin
        d11ctime_counter <= (d11ctime_counter - 1'd1);
    end
    if (susres_soft_int_clear) begin
        susres_soft_int_pending <= 1'd0;
    end
    susres_soft_int_trigger_d <= susres_soft_int_trigger;
    if (((~susres_soft_int_trigger) & susres_soft_int_trigger_d)) begin
        susres_soft_int_pending <= 1'd1;
    end
    if (always_on_rst) begin
        cpu_int_active <= 1'd0;
        irqarray0_eventsourceflex0_pending <= 1'd0;
        irqarray0_eventsourceflex0_trigger_d <= 1'd0;
        irqarray0_eventsourceflex1_pending <= 1'd0;
        irqarray0_eventsourceflex1_trigger_d <= 1'd0;
        irqarray0_eventsourceflex2_pending <= 1'd0;
        irqarray0_eventsourceflex2_trigger_d <= 1'd0;
        irqarray0_eventsourceflex3_pending <= 1'd0;
        irqarray0_eventsourceflex3_trigger_d <= 1'd0;
        irqarray0_eventsourceflex4_pending <= 1'd0;
        irqarray0_eventsourceflex4_trigger_d <= 1'd0;
        irqarray0_eventsourceflex5_pending <= 1'd0;
        irqarray0_eventsourceflex5_trigger_d <= 1'd0;
        irqarray0_eventsourceflex6_pending <= 1'd0;
        irqarray0_eventsourceflex6_trigger_d <= 1'd0;
        irqarray0_eventsourceflex7_pending <= 1'd0;
        irqarray0_eventsourceflex7_trigger_d <= 1'd0;
        irqarray0_eventsourceflex8_pending <= 1'd0;
        irqarray0_eventsourceflex8_trigger_d <= 1'd0;
        irqarray0_eventsourceflex9_pending <= 1'd0;
        irqarray0_eventsourceflex9_trigger_d <= 1'd0;
        irqarray0_eventsourceflex10_pending <= 1'd0;
        irqarray0_eventsourceflex10_trigger_d <= 1'd0;
        irqarray0_eventsourceflex11_pending <= 1'd0;
        irqarray0_eventsourceflex11_trigger_d <= 1'd0;
        irqarray0_eventsourceflex12_pending <= 1'd0;
        irqarray0_eventsourceflex12_trigger_d <= 1'd0;
        irqarray0_eventsourceflex13_pending <= 1'd0;
        irqarray0_eventsourceflex13_trigger_d <= 1'd0;
        irqarray0_eventsourceflex14_pending <= 1'd0;
        irqarray0_eventsourceflex14_trigger_d <= 1'd0;
        irqarray0_eventsourceflex15_pending <= 1'd0;
        irqarray0_eventsourceflex15_trigger_d <= 1'd0;
        irqarray1_eventsourceflex16_pending <= 1'd0;
        irqarray1_eventsourceflex16_trigger_d <= 1'd0;
        irqarray1_eventsourceflex17_pending <= 1'd0;
        irqarray1_eventsourceflex17_trigger_d <= 1'd0;
        irqarray1_eventsourceflex18_pending <= 1'd0;
        irqarray1_eventsourceflex18_trigger_d <= 1'd0;
        irqarray1_eventsourceflex19_pending <= 1'd0;
        irqarray1_eventsourceflex19_trigger_d <= 1'd0;
        irqarray1_eventsourceflex20_pending <= 1'd0;
        irqarray1_eventsourceflex20_trigger_d <= 1'd0;
        irqarray1_eventsourceflex21_pending <= 1'd0;
        irqarray1_eventsourceflex21_trigger_d <= 1'd0;
        irqarray1_eventsourceflex22_pending <= 1'd0;
        irqarray1_eventsourceflex22_trigger_d <= 1'd0;
        irqarray1_eventsourceflex23_pending <= 1'd0;
        irqarray1_eventsourceflex23_trigger_d <= 1'd0;
        irqarray1_eventsourceflex24_pending <= 1'd0;
        irqarray1_eventsourceflex24_trigger_d <= 1'd0;
        irqarray1_eventsourceflex25_pending <= 1'd0;
        irqarray1_eventsourceflex25_trigger_d <= 1'd0;
        irqarray1_eventsourceflex26_pending <= 1'd0;
        irqarray1_eventsourceflex26_trigger_d <= 1'd0;
        irqarray1_eventsourceflex27_pending <= 1'd0;
        irqarray1_eventsourceflex27_trigger_d <= 1'd0;
        irqarray1_eventsourceflex28_pending <= 1'd0;
        irqarray1_eventsourceflex28_trigger_d <= 1'd0;
        irqarray1_eventsourceflex29_pending <= 1'd0;
        irqarray1_eventsourceflex29_trigger_d <= 1'd0;
        irqarray1_eventsourceflex30_pending <= 1'd0;
        irqarray1_eventsourceflex30_trigger_d <= 1'd0;
        irqarray1_eventsourceflex31_pending <= 1'd0;
        irqarray1_eventsourceflex31_trigger_d <= 1'd0;
        irqarray2_eventsourceflex32_pending <= 1'd0;
        irqarray2_eventsourceflex32_trigger_d <= 1'd0;
        irqarray2_eventsourceflex33_pending <= 1'd0;
        irqarray2_eventsourceflex33_trigger_d <= 1'd0;
        irqarray2_eventsourceflex34_pending <= 1'd0;
        irqarray2_eventsourceflex34_trigger_d <= 1'd0;
        irqarray2_eventsourceflex35_pending <= 1'd0;
        irqarray2_eventsourceflex35_trigger_d <= 1'd0;
        irqarray2_eventsourceflex36_pending <= 1'd0;
        irqarray2_eventsourceflex36_trigger_d <= 1'd0;
        irqarray2_eventsourceflex37_pending <= 1'd0;
        irqarray2_eventsourceflex37_trigger_d <= 1'd0;
        irqarray2_eventsourceflex38_pending <= 1'd0;
        irqarray2_eventsourceflex38_trigger_d <= 1'd0;
        irqarray2_eventsourceflex39_pending <= 1'd0;
        irqarray2_eventsourceflex39_trigger_d <= 1'd0;
        irqarray2_eventsourceflex40_pending <= 1'd0;
        irqarray2_eventsourceflex40_trigger_d <= 1'd0;
        irqarray2_eventsourceflex41_pending <= 1'd0;
        irqarray2_eventsourceflex41_trigger_d <= 1'd0;
        irqarray2_eventsourceflex42_pending <= 1'd0;
        irqarray2_eventsourceflex42_trigger_d <= 1'd0;
        irqarray2_eventsourceflex43_pending <= 1'd0;
        irqarray2_eventsourceflex43_trigger_d <= 1'd0;
        irqarray2_eventsourceflex44_pending <= 1'd0;
        irqarray2_eventsourceflex44_trigger_d <= 1'd0;
        irqarray2_eventsourceflex45_pending <= 1'd0;
        irqarray2_eventsourceflex45_trigger_d <= 1'd0;
        irqarray2_eventsourceflex46_pending <= 1'd0;
        irqarray2_eventsourceflex46_trigger_d <= 1'd0;
        irqarray2_eventsourceflex47_pending <= 1'd0;
        irqarray2_eventsourceflex47_trigger_d <= 1'd0;
        irqarray3_eventsourceflex48_pending <= 1'd0;
        irqarray3_eventsourceflex48_trigger_d <= 1'd0;
        irqarray3_eventsourceflex49_pending <= 1'd0;
        irqarray3_eventsourceflex49_trigger_d <= 1'd0;
        irqarray3_eventsourceflex50_pending <= 1'd0;
        irqarray3_eventsourceflex50_trigger_d <= 1'd0;
        irqarray3_eventsourceflex51_pending <= 1'd0;
        irqarray3_eventsourceflex51_trigger_d <= 1'd0;
        irqarray3_eventsourceflex52_pending <= 1'd0;
        irqarray3_eventsourceflex52_trigger_d <= 1'd0;
        irqarray3_eventsourceflex53_pending <= 1'd0;
        irqarray3_eventsourceflex53_trigger_d <= 1'd0;
        irqarray3_eventsourceflex54_pending <= 1'd0;
        irqarray3_eventsourceflex54_trigger_d <= 1'd0;
        irqarray3_eventsourceflex55_pending <= 1'd0;
        irqarray3_eventsourceflex55_trigger_d <= 1'd0;
        irqarray3_eventsourceflex56_pending <= 1'd0;
        irqarray3_eventsourceflex56_trigger_d <= 1'd0;
        irqarray3_eventsourceflex57_pending <= 1'd0;
        irqarray3_eventsourceflex57_trigger_d <= 1'd0;
        irqarray3_eventsourceflex58_pending <= 1'd0;
        irqarray3_eventsourceflex58_trigger_d <= 1'd0;
        irqarray3_eventsourceflex59_pending <= 1'd0;
        irqarray3_eventsourceflex59_trigger_d <= 1'd0;
        irqarray3_eventsourceflex60_pending <= 1'd0;
        irqarray3_eventsourceflex60_trigger_d <= 1'd0;
        irqarray3_eventsourceflex61_pending <= 1'd0;
        irqarray3_eventsourceflex61_trigger_d <= 1'd0;
        irqarray3_eventsourceflex62_pending <= 1'd0;
        irqarray3_eventsourceflex62_trigger_d <= 1'd0;
        irqarray3_eventsourceflex63_pending <= 1'd0;
        irqarray3_eventsourceflex63_trigger_d <= 1'd0;
        irqarray4_eventsourceflex64_pending <= 1'd0;
        irqarray4_eventsourceflex64_trigger_d <= 1'd0;
        irqarray4_eventsourceflex65_pending <= 1'd0;
        irqarray4_eventsourceflex65_trigger_d <= 1'd0;
        irqarray4_eventsourceflex66_pending <= 1'd0;
        irqarray4_eventsourceflex66_trigger_d <= 1'd0;
        irqarray4_eventsourceflex67_pending <= 1'd0;
        irqarray4_eventsourceflex67_trigger_d <= 1'd0;
        irqarray4_eventsourceflex68_pending <= 1'd0;
        irqarray4_eventsourceflex68_trigger_d <= 1'd0;
        irqarray4_eventsourceflex69_pending <= 1'd0;
        irqarray4_eventsourceflex69_trigger_d <= 1'd0;
        irqarray4_eventsourceflex70_pending <= 1'd0;
        irqarray4_eventsourceflex70_trigger_d <= 1'd0;
        irqarray4_eventsourceflex71_pending <= 1'd0;
        irqarray4_eventsourceflex71_trigger_d <= 1'd0;
        irqarray4_eventsourceflex72_pending <= 1'd0;
        irqarray4_eventsourceflex72_trigger_d <= 1'd0;
        irqarray4_eventsourceflex73_pending <= 1'd0;
        irqarray4_eventsourceflex73_trigger_d <= 1'd0;
        irqarray4_eventsourceflex74_pending <= 1'd0;
        irqarray4_eventsourceflex74_trigger_d <= 1'd0;
        irqarray4_eventsourceflex75_pending <= 1'd0;
        irqarray4_eventsourceflex75_trigger_d <= 1'd0;
        irqarray4_eventsourceflex76_pending <= 1'd0;
        irqarray4_eventsourceflex76_trigger_d <= 1'd0;
        irqarray4_eventsourceflex77_pending <= 1'd0;
        irqarray4_eventsourceflex77_trigger_d <= 1'd0;
        irqarray4_eventsourceflex78_pending <= 1'd0;
        irqarray4_eventsourceflex78_trigger_d <= 1'd0;
        irqarray4_eventsourceflex79_pending <= 1'd0;
        irqarray4_eventsourceflex79_trigger_d <= 1'd0;
        irqarray5_eventsourceflex80_pending <= 1'd0;
        irqarray5_eventsourceflex80_trigger_d <= 1'd0;
        irqarray5_eventsourceflex81_pending <= 1'd0;
        irqarray5_eventsourceflex81_trigger_d <= 1'd0;
        irqarray5_eventsourceflex82_pending <= 1'd0;
        irqarray5_eventsourceflex82_trigger_d <= 1'd0;
        irqarray5_eventsourceflex83_pending <= 1'd0;
        irqarray5_eventsourceflex83_trigger_d <= 1'd0;
        irqarray5_eventsourceflex84_pending <= 1'd0;
        irqarray5_eventsourceflex84_trigger_d <= 1'd0;
        irqarray5_eventsourceflex85_pending <= 1'd0;
        irqarray5_eventsourceflex85_trigger_d <= 1'd0;
        irqarray5_eventsourceflex86_pending <= 1'd0;
        irqarray5_eventsourceflex86_trigger_d <= 1'd0;
        irqarray5_eventsourceflex87_pending <= 1'd0;
        irqarray5_eventsourceflex87_trigger_d <= 1'd0;
        irqarray5_eventsourceflex88_pending <= 1'd0;
        irqarray5_eventsourceflex88_trigger_d <= 1'd0;
        irqarray5_eventsourceflex89_pending <= 1'd0;
        irqarray5_eventsourceflex89_trigger_d <= 1'd0;
        irqarray5_eventsourceflex90_pending <= 1'd0;
        irqarray5_eventsourceflex90_trigger_d <= 1'd0;
        irqarray5_eventsourceflex91_pending <= 1'd0;
        irqarray5_eventsourceflex91_trigger_d <= 1'd0;
        irqarray5_eventsourceflex92_pending <= 1'd0;
        irqarray5_eventsourceflex92_trigger_d <= 1'd0;
        irqarray5_eventsourceflex93_pending <= 1'd0;
        irqarray5_eventsourceflex93_trigger_d <= 1'd0;
        irqarray5_eventsourceflex94_pending <= 1'd0;
        irqarray5_eventsourceflex94_trigger_d <= 1'd0;
        irqarray5_eventsourceflex95_pending <= 1'd0;
        irqarray5_eventsourceflex95_trigger_d <= 1'd0;
        irqarray6_eventsourceflex96_pending <= 1'd0;
        irqarray6_eventsourceflex96_trigger_d <= 1'd0;
        irqarray6_eventsourceflex97_pending <= 1'd0;
        irqarray6_eventsourceflex97_trigger_d <= 1'd0;
        irqarray6_eventsourceflex98_pending <= 1'd0;
        irqarray6_eventsourceflex98_trigger_d <= 1'd0;
        irqarray6_eventsourceflex99_pending <= 1'd0;
        irqarray6_eventsourceflex99_trigger_d <= 1'd0;
        irqarray6_eventsourceflex100_pending <= 1'd0;
        irqarray6_eventsourceflex100_trigger_d <= 1'd0;
        irqarray6_eventsourceflex101_pending <= 1'd0;
        irqarray6_eventsourceflex101_trigger_d <= 1'd0;
        irqarray6_eventsourceflex102_pending <= 1'd0;
        irqarray6_eventsourceflex102_trigger_d <= 1'd0;
        irqarray6_eventsourceflex103_pending <= 1'd0;
        irqarray6_eventsourceflex103_trigger_d <= 1'd0;
        irqarray6_eventsourceflex104_pending <= 1'd0;
        irqarray6_eventsourceflex104_trigger_d <= 1'd0;
        irqarray6_eventsourceflex105_pending <= 1'd0;
        irqarray6_eventsourceflex105_trigger_d <= 1'd0;
        irqarray6_eventsourceflex106_pending <= 1'd0;
        irqarray6_eventsourceflex106_trigger_d <= 1'd0;
        irqarray6_eventsourceflex107_pending <= 1'd0;
        irqarray6_eventsourceflex107_trigger_d <= 1'd0;
        irqarray6_eventsourceflex108_pending <= 1'd0;
        irqarray6_eventsourceflex108_trigger_d <= 1'd0;
        irqarray6_eventsourceflex109_pending <= 1'd0;
        irqarray6_eventsourceflex109_trigger_d <= 1'd0;
        irqarray6_eventsourceflex110_pending <= 1'd0;
        irqarray6_eventsourceflex110_trigger_d <= 1'd0;
        irqarray6_eventsourceflex111_pending <= 1'd0;
        irqarray6_eventsourceflex111_trigger_d <= 1'd0;
        irqarray7_eventsourceflex112_pending <= 1'd0;
        irqarray7_eventsourceflex112_trigger_d <= 1'd0;
        irqarray7_eventsourceflex113_pending <= 1'd0;
        irqarray7_eventsourceflex113_trigger_d <= 1'd0;
        irqarray7_eventsourceflex114_pending <= 1'd0;
        irqarray7_eventsourceflex114_trigger_d <= 1'd0;
        irqarray7_eventsourceflex115_pending <= 1'd0;
        irqarray7_eventsourceflex115_trigger_d <= 1'd0;
        irqarray7_eventsourceflex116_pending <= 1'd0;
        irqarray7_eventsourceflex116_trigger_d <= 1'd0;
        irqarray7_eventsourceflex117_pending <= 1'd0;
        irqarray7_eventsourceflex117_trigger_d <= 1'd0;
        irqarray7_eventsourceflex118_pending <= 1'd0;
        irqarray7_eventsourceflex118_trigger_d <= 1'd0;
        irqarray7_eventsourceflex119_pending <= 1'd0;
        irqarray7_eventsourceflex119_trigger_d <= 1'd0;
        irqarray7_eventsourceflex120_pending <= 1'd0;
        irqarray7_eventsourceflex120_trigger_d <= 1'd0;
        irqarray7_eventsourceflex121_pending <= 1'd0;
        irqarray7_eventsourceflex121_trigger_d <= 1'd0;
        irqarray7_eventsourceflex122_pending <= 1'd0;
        irqarray7_eventsourceflex122_trigger_d <= 1'd0;
        irqarray7_eventsourceflex123_pending <= 1'd0;
        irqarray7_eventsourceflex123_trigger_d <= 1'd0;
        irqarray7_eventsourceflex124_pending <= 1'd0;
        irqarray7_eventsourceflex124_trigger_d <= 1'd0;
        irqarray7_eventsourceflex125_pending <= 1'd0;
        irqarray7_eventsourceflex125_trigger_d <= 1'd0;
        irqarray7_eventsourceflex126_pending <= 1'd0;
        irqarray7_eventsourceflex126_trigger_d <= 1'd0;
        irqarray7_eventsourceflex127_pending <= 1'd0;
        irqarray7_eventsourceflex127_trigger_d <= 1'd0;
        irqarray8_eventsourceflex128_pending <= 1'd0;
        irqarray8_eventsourceflex128_trigger_d <= 1'd0;
        irqarray8_eventsourceflex129_pending <= 1'd0;
        irqarray8_eventsourceflex129_trigger_d <= 1'd0;
        irqarray8_eventsourceflex130_pending <= 1'd0;
        irqarray8_eventsourceflex130_trigger_d <= 1'd0;
        irqarray8_eventsourceflex131_pending <= 1'd0;
        irqarray8_eventsourceflex131_trigger_d <= 1'd0;
        irqarray8_eventsourceflex132_pending <= 1'd0;
        irqarray8_eventsourceflex132_trigger_d <= 1'd0;
        irqarray8_eventsourceflex133_pending <= 1'd0;
        irqarray8_eventsourceflex133_trigger_d <= 1'd0;
        irqarray8_eventsourceflex134_pending <= 1'd0;
        irqarray8_eventsourceflex134_trigger_d <= 1'd0;
        irqarray8_eventsourceflex135_pending <= 1'd0;
        irqarray8_eventsourceflex135_trigger_d <= 1'd0;
        irqarray8_eventsourceflex136_pending <= 1'd0;
        irqarray8_eventsourceflex136_trigger_d <= 1'd0;
        irqarray8_eventsourceflex137_pending <= 1'd0;
        irqarray8_eventsourceflex137_trigger_d <= 1'd0;
        irqarray8_eventsourceflex138_pending <= 1'd0;
        irqarray8_eventsourceflex138_trigger_d <= 1'd0;
        irqarray8_eventsourceflex139_pending <= 1'd0;
        irqarray8_eventsourceflex139_trigger_d <= 1'd0;
        irqarray8_eventsourceflex140_pending <= 1'd0;
        irqarray8_eventsourceflex140_trigger_d <= 1'd0;
        irqarray8_eventsourceflex141_pending <= 1'd0;
        irqarray8_eventsourceflex141_trigger_d <= 1'd0;
        irqarray8_eventsourceflex142_pending <= 1'd0;
        irqarray8_eventsourceflex142_trigger_d <= 1'd0;
        irqarray8_eventsourceflex143_pending <= 1'd0;
        irqarray8_eventsourceflex143_trigger_d <= 1'd0;
        irqarray9_eventsourceflex144_pending <= 1'd0;
        irqarray9_eventsourceflex144_trigger_d <= 1'd0;
        irqarray9_eventsourceflex145_pending <= 1'd0;
        irqarray9_eventsourceflex145_trigger_d <= 1'd0;
        irqarray9_eventsourceflex146_pending <= 1'd0;
        irqarray9_eventsourceflex146_trigger_d <= 1'd0;
        irqarray9_eventsourceflex147_pending <= 1'd0;
        irqarray9_eventsourceflex147_trigger_d <= 1'd0;
        irqarray9_eventsourceflex148_pending <= 1'd0;
        irqarray9_eventsourceflex148_trigger_d <= 1'd0;
        irqarray9_eventsourceflex149_pending <= 1'd0;
        irqarray9_eventsourceflex149_trigger_d <= 1'd0;
        irqarray9_eventsourceflex150_pending <= 1'd0;
        irqarray9_eventsourceflex150_trigger_d <= 1'd0;
        irqarray9_eventsourceflex151_pending <= 1'd0;
        irqarray9_eventsourceflex151_trigger_d <= 1'd0;
        irqarray9_eventsourceflex152_pending <= 1'd0;
        irqarray9_eventsourceflex152_trigger_d <= 1'd0;
        irqarray9_eventsourceflex153_pending <= 1'd0;
        irqarray9_eventsourceflex153_trigger_d <= 1'd0;
        irqarray9_eventsourceflex154_pending <= 1'd0;
        irqarray9_eventsourceflex154_trigger_d <= 1'd0;
        irqarray9_eventsourceflex155_pending <= 1'd0;
        irqarray9_eventsourceflex155_trigger_d <= 1'd0;
        irqarray9_eventsourceflex156_pending <= 1'd0;
        irqarray9_eventsourceflex156_trigger_d <= 1'd0;
        irqarray9_eventsourceflex157_pending <= 1'd0;
        irqarray9_eventsourceflex157_trigger_d <= 1'd0;
        irqarray9_eventsourceflex158_pending <= 1'd0;
        irqarray9_eventsourceflex158_trigger_d <= 1'd0;
        irqarray9_eventsourceflex159_pending <= 1'd0;
        irqarray9_eventsourceflex159_trigger_d <= 1'd0;
        irqarray10_eventsourceflex160_pending <= 1'd0;
        irqarray10_eventsourceflex160_trigger_d <= 1'd0;
        irqarray10_eventsourceflex161_pending <= 1'd0;
        irqarray10_eventsourceflex161_trigger_d <= 1'd0;
        irqarray10_eventsourceflex162_pending <= 1'd0;
        irqarray10_eventsourceflex162_trigger_d <= 1'd0;
        irqarray10_eventsourceflex163_pending <= 1'd0;
        irqarray10_eventsourceflex163_trigger_d <= 1'd0;
        irqarray10_eventsourceflex164_pending <= 1'd0;
        irqarray10_eventsourceflex164_trigger_d <= 1'd0;
        irqarray10_eventsourceflex165_pending <= 1'd0;
        irqarray10_eventsourceflex165_trigger_d <= 1'd0;
        irqarray10_eventsourceflex166_pending <= 1'd0;
        irqarray10_eventsourceflex166_trigger_d <= 1'd0;
        irqarray10_eventsourceflex167_pending <= 1'd0;
        irqarray10_eventsourceflex167_trigger_d <= 1'd0;
        irqarray10_eventsourceflex168_pending <= 1'd0;
        irqarray10_eventsourceflex168_trigger_d <= 1'd0;
        irqarray10_eventsourceflex169_pending <= 1'd0;
        irqarray10_eventsourceflex169_trigger_d <= 1'd0;
        irqarray10_eventsourceflex170_pending <= 1'd0;
        irqarray10_eventsourceflex170_trigger_d <= 1'd0;
        irqarray10_eventsourceflex171_pending <= 1'd0;
        irqarray10_eventsourceflex171_trigger_d <= 1'd0;
        irqarray10_eventsourceflex172_pending <= 1'd0;
        irqarray10_eventsourceflex172_trigger_d <= 1'd0;
        irqarray10_eventsourceflex173_pending <= 1'd0;
        irqarray10_eventsourceflex173_trigger_d <= 1'd0;
        irqarray10_eventsourceflex174_pending <= 1'd0;
        irqarray10_eventsourceflex174_trigger_d <= 1'd0;
        irqarray10_eventsourceflex175_pending <= 1'd0;
        irqarray10_eventsourceflex175_trigger_d <= 1'd0;
        irqarray11_eventsourceflex176_pending <= 1'd0;
        irqarray11_eventsourceflex176_trigger_d <= 1'd0;
        irqarray11_eventsourceflex177_pending <= 1'd0;
        irqarray11_eventsourceflex177_trigger_d <= 1'd0;
        irqarray11_eventsourceflex178_pending <= 1'd0;
        irqarray11_eventsourceflex178_trigger_d <= 1'd0;
        irqarray11_eventsourceflex179_pending <= 1'd0;
        irqarray11_eventsourceflex179_trigger_d <= 1'd0;
        irqarray11_eventsourceflex180_pending <= 1'd0;
        irqarray11_eventsourceflex180_trigger_d <= 1'd0;
        irqarray11_eventsourceflex181_pending <= 1'd0;
        irqarray11_eventsourceflex181_trigger_d <= 1'd0;
        irqarray11_eventsourceflex182_pending <= 1'd0;
        irqarray11_eventsourceflex182_trigger_d <= 1'd0;
        irqarray11_eventsourceflex183_pending <= 1'd0;
        irqarray11_eventsourceflex183_trigger_d <= 1'd0;
        irqarray11_eventsourceflex184_pending <= 1'd0;
        irqarray11_eventsourceflex184_trigger_d <= 1'd0;
        irqarray11_eventsourceflex185_pending <= 1'd0;
        irqarray11_eventsourceflex185_trigger_d <= 1'd0;
        irqarray11_eventsourceflex186_pending <= 1'd0;
        irqarray11_eventsourceflex186_trigger_d <= 1'd0;
        irqarray11_eventsourceflex187_pending <= 1'd0;
        irqarray11_eventsourceflex187_trigger_d <= 1'd0;
        irqarray11_eventsourceflex188_pending <= 1'd0;
        irqarray11_eventsourceflex188_trigger_d <= 1'd0;
        irqarray11_eventsourceflex189_pending <= 1'd0;
        irqarray11_eventsourceflex189_trigger_d <= 1'd0;
        irqarray11_eventsourceflex190_pending <= 1'd0;
        irqarray11_eventsourceflex190_trigger_d <= 1'd0;
        irqarray11_eventsourceflex191_pending <= 1'd0;
        irqarray11_eventsourceflex191_trigger_d <= 1'd0;
        irqarray12_eventsourceflex192_pending <= 1'd0;
        irqarray12_eventsourceflex192_trigger_d <= 1'd0;
        irqarray12_eventsourceflex193_pending <= 1'd0;
        irqarray12_eventsourceflex193_trigger_d <= 1'd0;
        irqarray12_eventsourceflex194_pending <= 1'd0;
        irqarray12_eventsourceflex194_trigger_d <= 1'd0;
        irqarray12_eventsourceflex195_pending <= 1'd0;
        irqarray12_eventsourceflex195_trigger_d <= 1'd0;
        irqarray12_eventsourceflex196_pending <= 1'd0;
        irqarray12_eventsourceflex196_trigger_d <= 1'd0;
        irqarray12_eventsourceflex197_pending <= 1'd0;
        irqarray12_eventsourceflex197_trigger_d <= 1'd0;
        irqarray12_eventsourceflex198_pending <= 1'd0;
        irqarray12_eventsourceflex198_trigger_d <= 1'd0;
        irqarray12_eventsourceflex199_pending <= 1'd0;
        irqarray12_eventsourceflex199_trigger_d <= 1'd0;
        irqarray12_eventsourceflex200_pending <= 1'd0;
        irqarray12_eventsourceflex200_trigger_d <= 1'd0;
        irqarray12_eventsourceflex201_pending <= 1'd0;
        irqarray12_eventsourceflex201_trigger_d <= 1'd0;
        irqarray12_eventsourceflex202_pending <= 1'd0;
        irqarray12_eventsourceflex202_trigger_d <= 1'd0;
        irqarray12_eventsourceflex203_pending <= 1'd0;
        irqarray12_eventsourceflex203_trigger_d <= 1'd0;
        irqarray12_eventsourceflex204_pending <= 1'd0;
        irqarray12_eventsourceflex204_trigger_d <= 1'd0;
        irqarray12_eventsourceflex205_pending <= 1'd0;
        irqarray12_eventsourceflex205_trigger_d <= 1'd0;
        irqarray12_eventsourceflex206_pending <= 1'd0;
        irqarray12_eventsourceflex206_trigger_d <= 1'd0;
        irqarray12_eventsourceflex207_pending <= 1'd0;
        irqarray12_eventsourceflex207_trigger_d <= 1'd0;
        irqarray13_eventsourceflex208_pending <= 1'd0;
        irqarray13_eventsourceflex208_trigger_d <= 1'd0;
        irqarray13_eventsourceflex209_pending <= 1'd0;
        irqarray13_eventsourceflex209_trigger_d <= 1'd0;
        irqarray13_eventsourceflex210_pending <= 1'd0;
        irqarray13_eventsourceflex210_trigger_d <= 1'd0;
        irqarray13_eventsourceflex211_pending <= 1'd0;
        irqarray13_eventsourceflex211_trigger_d <= 1'd0;
        irqarray13_eventsourceflex212_pending <= 1'd0;
        irqarray13_eventsourceflex212_trigger_d <= 1'd0;
        irqarray13_eventsourceflex213_pending <= 1'd0;
        irqarray13_eventsourceflex213_trigger_d <= 1'd0;
        irqarray13_eventsourceflex214_pending <= 1'd0;
        irqarray13_eventsourceflex214_trigger_d <= 1'd0;
        irqarray13_eventsourceflex215_pending <= 1'd0;
        irqarray13_eventsourceflex215_trigger_d <= 1'd0;
        irqarray13_eventsourceflex216_pending <= 1'd0;
        irqarray13_eventsourceflex216_trigger_d <= 1'd0;
        irqarray13_eventsourceflex217_pending <= 1'd0;
        irqarray13_eventsourceflex217_trigger_d <= 1'd0;
        irqarray13_eventsourceflex218_pending <= 1'd0;
        irqarray13_eventsourceflex218_trigger_d <= 1'd0;
        irqarray13_eventsourceflex219_pending <= 1'd0;
        irqarray13_eventsourceflex219_trigger_d <= 1'd0;
        irqarray13_eventsourceflex220_pending <= 1'd0;
        irqarray13_eventsourceflex220_trigger_d <= 1'd0;
        irqarray13_eventsourceflex221_pending <= 1'd0;
        irqarray13_eventsourceflex221_trigger_d <= 1'd0;
        irqarray13_eventsourceflex222_pending <= 1'd0;
        irqarray13_eventsourceflex222_trigger_d <= 1'd0;
        irqarray13_eventsourceflex223_pending <= 1'd0;
        irqarray13_eventsourceflex223_trigger_d <= 1'd0;
        irqarray14_eventsourceflex224_pending <= 1'd0;
        irqarray14_eventsourceflex224_trigger_d <= 1'd0;
        irqarray14_eventsourceflex225_pending <= 1'd0;
        irqarray14_eventsourceflex225_trigger_d <= 1'd0;
        irqarray14_eventsourceflex226_pending <= 1'd0;
        irqarray14_eventsourceflex226_trigger_d <= 1'd0;
        irqarray14_eventsourceflex227_pending <= 1'd0;
        irqarray14_eventsourceflex227_trigger_d <= 1'd0;
        irqarray14_eventsourceflex228_pending <= 1'd0;
        irqarray14_eventsourceflex228_trigger_d <= 1'd0;
        irqarray14_eventsourceflex229_pending <= 1'd0;
        irqarray14_eventsourceflex229_trigger_d <= 1'd0;
        irqarray14_eventsourceflex230_pending <= 1'd0;
        irqarray14_eventsourceflex230_trigger_d <= 1'd0;
        irqarray14_eventsourceflex231_pending <= 1'd0;
        irqarray14_eventsourceflex231_trigger_d <= 1'd0;
        irqarray14_eventsourceflex232_pending <= 1'd0;
        irqarray14_eventsourceflex232_trigger_d <= 1'd0;
        irqarray14_eventsourceflex233_pending <= 1'd0;
        irqarray14_eventsourceflex233_trigger_d <= 1'd0;
        irqarray14_eventsourceflex234_pending <= 1'd0;
        irqarray14_eventsourceflex234_trigger_d <= 1'd0;
        irqarray14_eventsourceflex235_pending <= 1'd0;
        irqarray14_eventsourceflex235_trigger_d <= 1'd0;
        irqarray14_eventsourceflex236_pending <= 1'd0;
        irqarray14_eventsourceflex236_trigger_d <= 1'd0;
        irqarray14_eventsourceflex237_pending <= 1'd0;
        irqarray14_eventsourceflex237_trigger_d <= 1'd0;
        irqarray14_eventsourceflex238_pending <= 1'd0;
        irqarray14_eventsourceflex238_trigger_d <= 1'd0;
        irqarray14_eventsourceflex239_pending <= 1'd0;
        irqarray14_eventsourceflex239_trigger_d <= 1'd0;
        irqarray15_eventsourceflex240_pending <= 1'd0;
        irqarray15_eventsourceflex240_trigger_d <= 1'd0;
        irqarray15_eventsourceflex241_pending <= 1'd0;
        irqarray15_eventsourceflex241_trigger_d <= 1'd0;
        irqarray15_eventsourceflex242_pending <= 1'd0;
        irqarray15_eventsourceflex242_trigger_d <= 1'd0;
        irqarray15_eventsourceflex243_pending <= 1'd0;
        irqarray15_eventsourceflex243_trigger_d <= 1'd0;
        irqarray15_eventsourceflex244_pending <= 1'd0;
        irqarray15_eventsourceflex244_trigger_d <= 1'd0;
        irqarray15_eventsourceflex245_pending <= 1'd0;
        irqarray15_eventsourceflex245_trigger_d <= 1'd0;
        irqarray15_eventsourceflex246_pending <= 1'd0;
        irqarray15_eventsourceflex246_trigger_d <= 1'd0;
        irqarray15_eventsourceflex247_pending <= 1'd0;
        irqarray15_eventsourceflex247_trigger_d <= 1'd0;
        irqarray15_eventsourceflex248_pending <= 1'd0;
        irqarray15_eventsourceflex248_trigger_d <= 1'd0;
        irqarray15_eventsourceflex249_pending <= 1'd0;
        irqarray15_eventsourceflex249_trigger_d <= 1'd0;
        irqarray15_eventsourceflex250_pending <= 1'd0;
        irqarray15_eventsourceflex250_trigger_d <= 1'd0;
        irqarray15_eventsourceflex251_pending <= 1'd0;
        irqarray15_eventsourceflex251_trigger_d <= 1'd0;
        irqarray15_eventsourceflex252_pending <= 1'd0;
        irqarray15_eventsourceflex252_trigger_d <= 1'd0;
        irqarray15_eventsourceflex253_pending <= 1'd0;
        irqarray15_eventsourceflex253_trigger_d <= 1'd0;
        irqarray15_eventsourceflex254_pending <= 1'd0;
        irqarray15_eventsourceflex254_trigger_d <= 1'd0;
        irqarray15_eventsourceflex255_pending <= 1'd0;
        irqarray15_eventsourceflex255_trigger_d <= 1'd0;
        irqarray16_eventsourceflex256_pending <= 1'd0;
        irqarray16_eventsourceflex256_trigger_d <= 1'd0;
        irqarray16_eventsourceflex257_pending <= 1'd0;
        irqarray16_eventsourceflex257_trigger_d <= 1'd0;
        irqarray16_eventsourceflex258_pending <= 1'd0;
        irqarray16_eventsourceflex258_trigger_d <= 1'd0;
        irqarray16_eventsourceflex259_pending <= 1'd0;
        irqarray16_eventsourceflex259_trigger_d <= 1'd0;
        irqarray16_eventsourceflex260_pending <= 1'd0;
        irqarray16_eventsourceflex260_trigger_d <= 1'd0;
        irqarray16_eventsourceflex261_pending <= 1'd0;
        irqarray16_eventsourceflex261_trigger_d <= 1'd0;
        irqarray16_eventsourceflex262_pending <= 1'd0;
        irqarray16_eventsourceflex262_trigger_d <= 1'd0;
        irqarray16_eventsourceflex263_pending <= 1'd0;
        irqarray16_eventsourceflex263_trigger_d <= 1'd0;
        irqarray16_eventsourceflex264_pending <= 1'd0;
        irqarray16_eventsourceflex264_trigger_d <= 1'd0;
        irqarray16_eventsourceflex265_pending <= 1'd0;
        irqarray16_eventsourceflex265_trigger_d <= 1'd0;
        irqarray16_eventsourceflex266_pending <= 1'd0;
        irqarray16_eventsourceflex266_trigger_d <= 1'd0;
        irqarray16_eventsourceflex267_pending <= 1'd0;
        irqarray16_eventsourceflex267_trigger_d <= 1'd0;
        irqarray16_eventsourceflex268_pending <= 1'd0;
        irqarray16_eventsourceflex268_trigger_d <= 1'd0;
        irqarray16_eventsourceflex269_pending <= 1'd0;
        irqarray16_eventsourceflex269_trigger_d <= 1'd0;
        irqarray16_eventsourceflex270_pending <= 1'd0;
        irqarray16_eventsourceflex270_trigger_d <= 1'd0;
        irqarray16_eventsourceflex271_pending <= 1'd0;
        irqarray16_eventsourceflex271_trigger_d <= 1'd0;
        irqarray17_eventsourceflex272_pending <= 1'd0;
        irqarray17_eventsourceflex272_trigger_d <= 1'd0;
        irqarray17_eventsourceflex273_pending <= 1'd0;
        irqarray17_eventsourceflex273_trigger_d <= 1'd0;
        irqarray17_eventsourceflex274_pending <= 1'd0;
        irqarray17_eventsourceflex274_trigger_d <= 1'd0;
        irqarray17_eventsourceflex275_pending <= 1'd0;
        irqarray17_eventsourceflex275_trigger_d <= 1'd0;
        irqarray17_eventsourceflex276_pending <= 1'd0;
        irqarray17_eventsourceflex276_trigger_d <= 1'd0;
        irqarray17_eventsourceflex277_pending <= 1'd0;
        irqarray17_eventsourceflex277_trigger_d <= 1'd0;
        irqarray17_eventsourceflex278_pending <= 1'd0;
        irqarray17_eventsourceflex278_trigger_d <= 1'd0;
        irqarray17_eventsourceflex279_pending <= 1'd0;
        irqarray17_eventsourceflex279_trigger_d <= 1'd0;
        irqarray17_eventsourceflex280_pending <= 1'd0;
        irqarray17_eventsourceflex280_trigger_d <= 1'd0;
        irqarray17_eventsourceflex281_pending <= 1'd0;
        irqarray17_eventsourceflex281_trigger_d <= 1'd0;
        irqarray17_eventsourceflex282_pending <= 1'd0;
        irqarray17_eventsourceflex282_trigger_d <= 1'd0;
        irqarray17_eventsourceflex283_pending <= 1'd0;
        irqarray17_eventsourceflex283_trigger_d <= 1'd0;
        irqarray17_eventsourceflex284_pending <= 1'd0;
        irqarray17_eventsourceflex284_trigger_d <= 1'd0;
        irqarray17_eventsourceflex285_pending <= 1'd0;
        irqarray17_eventsourceflex285_trigger_d <= 1'd0;
        irqarray17_eventsourceflex286_pending <= 1'd0;
        irqarray17_eventsourceflex286_trigger_d <= 1'd0;
        irqarray17_eventsourceflex287_pending <= 1'd0;
        irqarray17_eventsourceflex287_trigger_d <= 1'd0;
        irqarray18_eventsourceflex288_pending <= 1'd0;
        irqarray18_eventsourceflex288_trigger_d <= 1'd0;
        irqarray18_eventsourceflex289_pending <= 1'd0;
        irqarray18_eventsourceflex289_trigger_d <= 1'd0;
        irqarray18_eventsourceflex290_pending <= 1'd0;
        irqarray18_eventsourceflex290_trigger_d <= 1'd0;
        irqarray18_eventsourceflex291_pending <= 1'd0;
        irqarray18_eventsourceflex291_trigger_d <= 1'd0;
        irqarray18_eventsourceflex292_pending <= 1'd0;
        irqarray18_eventsourceflex292_trigger_d <= 1'd0;
        irqarray18_eventsourceflex293_pending <= 1'd0;
        irqarray18_eventsourceflex293_trigger_d <= 1'd0;
        irqarray18_eventsourceflex294_pending <= 1'd0;
        irqarray18_eventsourceflex294_trigger_d <= 1'd0;
        irqarray18_eventsourceflex295_pending <= 1'd0;
        irqarray18_eventsourceflex295_trigger_d <= 1'd0;
        irqarray18_eventsourceflex296_pending <= 1'd0;
        irqarray18_eventsourceflex296_trigger_d <= 1'd0;
        irqarray18_eventsourceflex297_pending <= 1'd0;
        irqarray18_eventsourceflex297_trigger_d <= 1'd0;
        irqarray18_eventsourceflex298_pending <= 1'd0;
        irqarray18_eventsourceflex298_trigger_d <= 1'd0;
        irqarray18_eventsourceflex299_pending <= 1'd0;
        irqarray18_eventsourceflex299_trigger_d <= 1'd0;
        irqarray18_eventsourceflex300_pending <= 1'd0;
        irqarray18_eventsourceflex300_trigger_d <= 1'd0;
        irqarray18_eventsourceflex301_pending <= 1'd0;
        irqarray18_eventsourceflex301_trigger_d <= 1'd0;
        irqarray18_eventsourceflex302_pending <= 1'd0;
        irqarray18_eventsourceflex302_trigger_d <= 1'd0;
        irqarray18_eventsourceflex303_pending <= 1'd0;
        irqarray18_eventsourceflex303_trigger_d <= 1'd0;
        irqarray19_eventsourceflex304_pending <= 1'd0;
        irqarray19_eventsourceflex304_trigger_d <= 1'd0;
        irqarray19_eventsourceflex305_pending <= 1'd0;
        irqarray19_eventsourceflex305_trigger_d <= 1'd0;
        irqarray19_eventsourceflex306_pending <= 1'd0;
        irqarray19_eventsourceflex306_trigger_d <= 1'd0;
        irqarray19_eventsourceflex307_pending <= 1'd0;
        irqarray19_eventsourceflex307_trigger_d <= 1'd0;
        irqarray19_eventsourceflex308_pending <= 1'd0;
        irqarray19_eventsourceflex308_trigger_d <= 1'd0;
        irqarray19_eventsourceflex309_pending <= 1'd0;
        irqarray19_eventsourceflex309_trigger_d <= 1'd0;
        irqarray19_eventsourceflex310_pending <= 1'd0;
        irqarray19_eventsourceflex310_trigger_d <= 1'd0;
        irqarray19_eventsourceflex311_pending <= 1'd0;
        irqarray19_eventsourceflex311_trigger_d <= 1'd0;
        irqarray19_eventsourceflex312_pending <= 1'd0;
        irqarray19_eventsourceflex312_trigger_d <= 1'd0;
        irqarray19_eventsourceflex313_pending <= 1'd0;
        irqarray19_eventsourceflex313_trigger_d <= 1'd0;
        irqarray19_eventsourceflex314_pending <= 1'd0;
        irqarray19_eventsourceflex314_trigger_d <= 1'd0;
        irqarray19_eventsourceflex315_pending <= 1'd0;
        irqarray19_eventsourceflex315_trigger_d <= 1'd0;
        irqarray19_eventsourceflex316_pending <= 1'd0;
        irqarray19_eventsourceflex316_trigger_d <= 1'd0;
        irqarray19_eventsourceflex317_pending <= 1'd0;
        irqarray19_eventsourceflex317_trigger_d <= 1'd0;
        irqarray19_eventsourceflex318_pending <= 1'd0;
        irqarray19_eventsourceflex318_trigger_d <= 1'd0;
        irqarray19_eventsourceflex319_pending <= 1'd0;
        irqarray19_eventsourceflex319_trigger_d <= 1'd0;
        ticktimer_prescaler <= 32'd800000;
        ticktimer_timer0 <= 64'd0;
        ticktimer_load_xfer_ps_toggle_i <= 1'd0;
        ticktimer_load_xfer_ps_ack_toggle_i <= 1'd0;
        ticktimer_load_xfer_blind <= 1'd0;
        ticktimer_paused1 <= 1'd0;
        ticktimer_timer_sync_starter <= 1'd1;
        ticktimer_timer_sync_ping_toggle_i <= 1'd0;
        ticktimer_timer_sync_ping_o1 <= 1'd0;
        ticktimer_timer_sync_pong_toggle_i <= 1'd0;
        ticktimer_timer_sync_count <= 8'd128;
        ticktimer_resume_sync_starter <= 1'd1;
        ticktimer_resume_sync_ping_toggle_i <= 1'd0;
        ticktimer_resume_sync_ping_o1 <= 1'd0;
        ticktimer_resume_sync_pong_toggle_i <= 1'd0;
        ticktimer_resume_sync_count <= 8'd128;
        ticktimer_reset_xfer_ps_toggle_i <= 1'd0;
        ticktimer_reset_xfer_ps_ack_toggle_i <= 1'd0;
        ticktimer_reset_xfer_blind <= 1'd0;
        ticktimer_ping_ps_toggle_i <= 1'd0;
        ticktimer_ping_ps_ack_toggle_i <= 1'd0;
        ticktimer_ping_blind <= 1'd0;
        ticktimer_pong_ps_toggle_i <= 1'd0;
        ticktimer_pong_ps_ack_toggle_i <= 1'd0;
        ticktimer_pong_blind <= 1'd0;
        ticktimer_lockout_alarm <= 1'd0;
        ticktimer_alarm3 <= 1'd0;
        ticktimer_target_xfer_starter <= 1'd1;
        ticktimer_target_xfer_ping_toggle_i <= 1'd0;
        ticktimer_target_xfer_ping_o1 <= 1'd0;
        ticktimer_target_xfer_pong_toggle_i <= 1'd0;
        ticktimer_target_xfer_count <= 8'd128;
        d11ctime_counter <= 32'd400000;
        d11ctime_heartbeat <= 1'd0;
        susres_soft_int_pending <= 1'd0;
        susres_soft_int_trigger_d <= 1'd0;
    end
    multiregimpl0_regs0 <= ticktimer_pause0;
    multiregimpl0_regs1 <= multiregimpl0_regs0;
    multiregimpl1_regs0 <= ticktimer_load_xfer_ps_toggle_i;
    multiregimpl1_regs1 <= multiregimpl1_regs0;
    multiregimpl2_regs0 <= ticktimer_load_xfer_ps_ack_toggle_i;
    multiregimpl2_regs1 <= multiregimpl2_regs0;
    multiregimpl3_regs0 <= ticktimer_paused1;
    multiregimpl3_regs1 <= multiregimpl3_regs0;
    multiregimpl4_regs0 <= ticktimer_timer_sync_ping_toggle_i;
    multiregimpl4_regs1 <= multiregimpl4_regs0;
    multiregimpl5_regs0 <= ticktimer_timer_sync_pong_toggle_i;
    multiregimpl5_regs1 <= multiregimpl5_regs0;
    multiregimpl6_regs0 <= ticktimer_timer_sync_ibuffer;
    multiregimpl6_regs1 <= multiregimpl6_regs0;
    multiregimpl7_regs0 <= ticktimer_resume_sync_ping_toggle_i;
    multiregimpl7_regs1 <= multiregimpl7_regs0;
    multiregimpl8_regs0 <= ticktimer_resume_sync_pong_toggle_i;
    multiregimpl8_regs1 <= multiregimpl8_regs0;
    multiregimpl9_regs0 <= ticktimer_resume_sync_ibuffer;
    multiregimpl9_regs1 <= multiregimpl9_regs0;
    multiregimpl10_regs0 <= ticktimer_reset_xfer_ps_toggle_i;
    multiregimpl10_regs1 <= multiregimpl10_regs0;
    multiregimpl11_regs0 <= ticktimer_reset_xfer_ps_ack_toggle_i;
    multiregimpl11_regs1 <= multiregimpl11_regs0;
    multiregimpl12_regs0 <= ticktimer_ping_ps_toggle_i;
    multiregimpl12_regs1 <= multiregimpl12_regs0;
    multiregimpl13_regs0 <= ticktimer_ping_ps_ack_toggle_i;
    multiregimpl13_regs1 <= multiregimpl13_regs0;
    multiregimpl14_regs0 <= ticktimer_pong_ps_toggle_i;
    multiregimpl14_regs1 <= multiregimpl14_regs0;
    multiregimpl15_regs0 <= ticktimer_pong_ps_ack_toggle_i;
    multiregimpl15_regs1 <= multiregimpl15_regs0;
    multiregimpl16_regs0 <= ticktimer_target_xfer_ping_toggle_i;
    multiregimpl16_regs1 <= multiregimpl16_regs0;
    multiregimpl17_regs0 <= ticktimer_target_xfer_pong_toggle_i;
    multiregimpl17_regs1 <= multiregimpl17_regs0;
    multiregimpl18_regs0 <= ticktimer_target_xfer_ibuffer;
    multiregimpl18_regs1 <= multiregimpl18_regs0;
end

always @(posedge sys_clk) begin
    if (cramsoc_ibus_axi_ar_valid) begin
        ibus_r_active <= 1'd1;
    end else begin
        if (((cramsoc_ibus_axi_r_valid & cramsoc_ibus_axi_r_ready) & cramsoc_ibus_axi_r_last)) begin
            ibus_r_active <= 1'd0;
        end
    end
    if (cramsoc_dbus_ar_valid) begin
        dbus_r_active <= 1'd1;
    end else begin
        if (((cramsoc_dbus_r_valid & cramsoc_dbus_r_ready) & cramsoc_dbus_r_last)) begin
            dbus_r_active <= 1'd0;
        end
    end
    if (cramsoc_dbus_aw_valid) begin
        dbus_w_active <= 1'd1;
    end else begin
        if ((cramsoc_dbus_b_valid & cramsoc_dbus_b_ready)) begin
            dbus_w_active <= 1'd0;
        end
    end
    if (cramsoc_peripherals_ar_valid) begin
        pbus_r_active <= 1'd1;
    end else begin
        if ((cramsoc_peripherals_r_valid & cramsoc_peripherals_r_ready)) begin
            pbus_r_active <= 1'd0;
        end
    end
    if (cramsoc_peripherals_aw_valid) begin
        pbus_w_active <= 1'd1;
    end else begin
        if ((cramsoc_peripherals_b_valid & cramsoc_peripherals_b_ready)) begin
            pbus_w_active <= 1'd0;
        end
    end
    if (axi_active) begin
        active_timeout <= 7'd64;
    end else begin
        if ((active_timeout > 1'd0)) begin
            active_timeout <= (active_timeout - 1'd1);
        end else begin
            active_timeout <= active_timeout;
        end
    end
    if (socbushandler_axiliterequestcounter0_empty) begin
        socbushandler_slave_sel_reg0 <= socbushandler_slave_sel_dec0;
    end
    if (socbushandler_axiliterequestcounter1_empty) begin
        socbushandler_slave_sel_reg1 <= socbushandler_slave_sel_dec1;
    end
    if (((cramsoc_corecsr_aw_valid & cramsoc_corecsr_aw_ready) & (cramsoc_corecsr_b_valid & cramsoc_corecsr_b_ready))) begin
        socbushandler_axiliterequestcounter0_counter <= socbushandler_axiliterequestcounter0_counter;
    end else begin
        if (((cramsoc_corecsr_aw_valid & cramsoc_corecsr_aw_ready) & (~socbushandler_axiliterequestcounter0_full))) begin
            socbushandler_axiliterequestcounter0_counter <= (socbushandler_axiliterequestcounter0_counter + 1'd1);
        end else begin
            if (((cramsoc_corecsr_b_valid & cramsoc_corecsr_b_ready) & (~socbushandler_axiliterequestcounter0_empty))) begin
                socbushandler_axiliterequestcounter0_counter <= (socbushandler_axiliterequestcounter0_counter - 1'd1);
            end
        end
    end
    if (((cramsoc_corecsr_ar_valid & cramsoc_corecsr_ar_ready) & (cramsoc_corecsr_r_valid & cramsoc_corecsr_r_ready))) begin
        socbushandler_axiliterequestcounter1_counter <= socbushandler_axiliterequestcounter1_counter;
    end else begin
        if (((cramsoc_corecsr_ar_valid & cramsoc_corecsr_ar_ready) & (~socbushandler_axiliterequestcounter1_full))) begin
            socbushandler_axiliterequestcounter1_counter <= (socbushandler_axiliterequestcounter1_counter + 1'd1);
        end else begin
            if (((cramsoc_corecsr_r_valid & cramsoc_corecsr_r_ready) & (~socbushandler_axiliterequestcounter1_empty))) begin
                socbushandler_axiliterequestcounter1_counter <= (socbushandler_axiliterequestcounter1_counter - 1'd1);
            end
        end
    end
    if (((cramsoc_aw_valid & cramsoc_aw_ready) & (cramsoc_b_valid & cramsoc_b_ready))) begin
        socbushandler_wr_lock_counter <= socbushandler_wr_lock_counter;
    end else begin
        if (((cramsoc_aw_valid & cramsoc_aw_ready) & (~socbushandler_wr_lock_full))) begin
            socbushandler_wr_lock_counter <= (socbushandler_wr_lock_counter + 1'd1);
        end else begin
            if (((cramsoc_b_valid & cramsoc_b_ready) & (~socbushandler_wr_lock_empty))) begin
                socbushandler_wr_lock_counter <= (socbushandler_wr_lock_counter - 1'd1);
            end
        end
    end
    if (((cramsoc_ar_valid & cramsoc_ar_ready) & (cramsoc_r_valid & cramsoc_r_ready))) begin
        socbushandler_rd_lock_counter <= socbushandler_rd_lock_counter;
    end else begin
        if (((cramsoc_ar_valid & cramsoc_ar_ready) & (~socbushandler_rd_lock_full))) begin
            socbushandler_rd_lock_counter <= (socbushandler_rd_lock_counter + 1'd1);
        end else begin
            if (((cramsoc_r_valid & cramsoc_r_ready) & (~socbushandler_rd_lock_empty))) begin
                socbushandler_rd_lock_counter <= (socbushandler_rd_lock_counter - 1'd1);
            end
        end
    end
    reset_debug_logic <= o_resetOut;
    debug_reset <= (reset_debug_logic | sys_rst);
    if (cramsoc_en_storage) begin
        if ((cramsoc_value == 1'd0)) begin
            cramsoc_value <= cramsoc_reload_storage;
        end else begin
            cramsoc_value <= (cramsoc_value - 1'd1);
        end
    end else begin
        cramsoc_value <= cramsoc_load_storage;
    end
    if (cramsoc_update_value_re) begin
        cramsoc_value_status <= cramsoc_value;
    end
    if (cramsoc_zero_clear) begin
        cramsoc_zero_pending <= 1'd0;
    end
    cramsoc_zero_trigger_d <= cramsoc_zero_trigger;
    if ((cramsoc_zero_trigger & (~cramsoc_zero_trigger_d))) begin
        cramsoc_zero_pending <= 1'd1;
    end
    if (sys_rst) begin
        if (trimming_reset_ena_1) begin
            latched_value <= trimming_reset_1;
        end else begin
            latched_value <= 31'd1610612736;
        end
    end else begin
        latched_value <= latched_value;
    end
    if (coreuser_protect) begin
        coreuser_enable1 <= coreuser_enable1;
        coreuser_invert_priv1 <= coreuser_invert_priv1;
        coreuser_lut01 <= coreuser_lut01;
        coreuser_lut11 <= coreuser_lut11;
        coreuser_lut21 <= coreuser_lut21;
        coreuser_lut31 <= coreuser_lut31;
        coreuser_lut41 <= coreuser_lut41;
        coreuser_lut51 <= coreuser_lut51;
        coreuser_lut61 <= coreuser_lut61;
        coreuser_lut71 <= coreuser_lut71;
        coreuser_user01 <= coreuser_user01;
        coreuser_user11 <= coreuser_user11;
        coreuser_user21 <= coreuser_user21;
        coreuser_user31 <= coreuser_user31;
        coreuser_user41 <= coreuser_user41;
        coreuser_user51 <= coreuser_user51;
        coreuser_user61 <= coreuser_user61;
        coreuser_user71 <= coreuser_user71;
        coreuser_user_default <= coreuser_user_default;
    end else begin
        coreuser_enable1 <= coreuser_enable0;
        coreuser_invert_priv1 <= coreuser_invert_priv0;
        coreuser_lut01 <= coreuser_lut00;
        coreuser_lut11 <= coreuser_lut10;
        coreuser_lut21 <= coreuser_lut20;
        coreuser_lut31 <= coreuser_lut30;
        coreuser_lut41 <= coreuser_lut40;
        coreuser_lut51 <= coreuser_lut50;
        coreuser_lut61 <= coreuser_lut60;
        coreuser_lut71 <= coreuser_lut70;
        coreuser_user01 <= coreuser_user00;
        coreuser_user11 <= coreuser_user10;
        coreuser_user21 <= coreuser_user20;
        coreuser_user31 <= coreuser_user30;
        coreuser_user41 <= coreuser_user40;
        coreuser_user51 <= coreuser_user50;
        coreuser_user61 <= coreuser_user60;
        coreuser_user71 <= coreuser_user70;
        coreuser_user_default <= coreuser_default;
    end
    coreuser_coreuser <= coreuser_vex;
    coreuser_mm <= vex_mm;
    coreuser_vex[7:4] <= coreuser_coreuser_4bit;
    coreuser_vex[3:0] <= {coreuser_coreuser_4bit[0], coreuser_coreuser_4bit[1], coreuser_coreuser_4bit[2], coreuser_coreuser_4bit[3]};
    if (coreuser_enable1) begin
        vex_mm <= ((cramsoc_privilege[0] | cramsoc_privilege[1]) ^ coreuser_invert_priv1);
    end else begin
        vex_mm <= default_mm;
    end
    if (mailbox_available_clear) begin
        mailbox_available_pending <= 1'd0;
    end
    if (mailbox_available_trigger) begin
        mailbox_available_pending <= 1'd1;
    end
    if (mailbox_abort_init_clear) begin
        mailbox_abort_init_pending <= 1'd0;
    end
    mailbox_abort_init_trigger_d <= mailbox_abort_init_trigger;
    if ((mailbox_abort_init_trigger & (~mailbox_abort_init_trigger_d))) begin
        mailbox_abort_init_pending <= 1'd1;
    end
    if (mailbox_abort_done_clear) begin
        mailbox_abort_done_pending <= 1'd0;
    end
    mailbox_abort_done_trigger_d <= mailbox_abort_done_trigger;
    if ((mailbox_abort_done_trigger & (~mailbox_abort_done_trigger_d))) begin
        mailbox_abort_done_pending <= 1'd1;
    end
    if (mailbox_error_clear) begin
        mailbox_error_pending <= 1'd0;
    end
    mailbox_error_trigger_d <= mailbox_error_trigger;
    if ((mailbox_error_trigger & (~mailbox_error_trigger_d))) begin
        mailbox_error_pending <= 1'd1;
    end
    if (mailbox_w_over_clear) begin
        mailbox_w_over_bit <= 1'd0;
    end else begin
        if (mailbox_w_over_flag) begin
            mailbox_w_over_bit <= 1'd1;
        end else begin
            mailbox_w_over_bit <= mailbox_w_over_bit;
        end
    end
    if (mailbox_syncfifobufferedmacro0_fifo_re) begin
        mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_readable <= 1'd1;
    end else begin
        if (mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_re) begin
            mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_readable <= 1'd0;
        end
    end
    if (($signed({1'd0, (mailbox_syncfifobufferedmacro0_fifo_we & mailbox_syncfifobufferedmacro0_fifo_writable)}) & -1'd1)) begin
        mailbox_syncfifobufferedmacro0_fifo_produce <= (mailbox_syncfifobufferedmacro0_fifo_produce + 1'd1);
    end
    if (mailbox_syncfifobufferedmacro0_fifo_do_read) begin
        mailbox_syncfifobufferedmacro0_fifo_consume <= (mailbox_syncfifobufferedmacro0_fifo_consume + 1'd1);
    end
    if (($signed({1'd0, (mailbox_syncfifobufferedmacro0_fifo_we & mailbox_syncfifobufferedmacro0_fifo_writable)}) & -1'd1)) begin
        if ((~mailbox_syncfifobufferedmacro0_fifo_do_read)) begin
            mailbox_syncfifobufferedmacro0_fifo_level <= (mailbox_syncfifobufferedmacro0_fifo_level + 1'd1);
        end
    end else begin
        if (mailbox_syncfifobufferedmacro0_fifo_do_read) begin
            mailbox_syncfifobufferedmacro0_fifo_level <= (mailbox_syncfifobufferedmacro0_fifo_level - 1'd1);
        end
    end
    if (mailbox_w_fifo_reset_sys) begin
        mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_readable <= 1'd0;
        mailbox_syncfifobufferedmacro0_fifo_level <= 11'd0;
        mailbox_syncfifobufferedmacro0_fifo_produce <= 10'd0;
        mailbox_syncfifobufferedmacro0_fifo_consume <= 10'd0;
    end
    if (mailbox_r_over_clear) begin
        mailbox_r_over_bit <= 1'd0;
    end else begin
        if (mailbox_r_over_flag) begin
            mailbox_r_over_bit <= 1'd1;
        end else begin
            mailbox_r_over_bit <= mailbox_r_over_bit;
        end
    end
    if (mailbox_syncfifobufferedmacro1_fifo_re) begin
        mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_readable <= 1'd1;
    end else begin
        if (mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_re) begin
            mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_readable <= 1'd0;
        end
    end
    if (($signed({1'd0, (mailbox_syncfifobufferedmacro1_fifo_we & mailbox_syncfifobufferedmacro1_fifo_writable)}) & -1'd1)) begin
        mailbox_syncfifobufferedmacro1_fifo_produce <= (mailbox_syncfifobufferedmacro1_fifo_produce + 1'd1);
    end
    if (mailbox_syncfifobufferedmacro1_fifo_do_read) begin
        mailbox_syncfifobufferedmacro1_fifo_consume <= (mailbox_syncfifobufferedmacro1_fifo_consume + 1'd1);
    end
    if (($signed({1'd0, (mailbox_syncfifobufferedmacro1_fifo_we & mailbox_syncfifobufferedmacro1_fifo_writable)}) & -1'd1)) begin
        if ((~mailbox_syncfifobufferedmacro1_fifo_do_read)) begin
            mailbox_syncfifobufferedmacro1_fifo_level <= (mailbox_syncfifobufferedmacro1_fifo_level + 1'd1);
        end
    end else begin
        if (mailbox_syncfifobufferedmacro1_fifo_do_read) begin
            mailbox_syncfifobufferedmacro1_fifo_level <= (mailbox_syncfifobufferedmacro1_fifo_level - 1'd1);
        end
    end
    if (mailbox_r_fifo_reset_sys) begin
        mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_readable <= 1'd0;
        mailbox_syncfifobufferedmacro1_fifo_level <= 11'd0;
        mailbox_syncfifobufferedmacro1_fifo_produce <= 10'd0;
        mailbox_syncfifobufferedmacro1_fifo_consume <= 10'd0;
    end
    cramsoc_mailbox_state <= cramsoc_mailbox_next_state;
    if (mailbox_abort_ack1_mailbox_next_value_ce0) begin
        mailbox_abort_ack1 <= mailbox_abort_ack1_mailbox_next_value0;
    end
    if (mailbox_abort_in_progress1_mailbox_next_value_ce1) begin
        mailbox_abort_in_progress1 <= mailbox_abort_in_progress1_mailbox_next_value1;
    end
    if (mailbox_w_abort_mailbox_next_value_ce2) begin
        mailbox_w_abort <= mailbox_w_abort_mailbox_next_value2;
    end
    if ((mb_client_wdata_re & (~mb_client_w_ready))) begin
        mb_client_w_pending <= 1'd1;
    end else begin
        if ((mb_client_w_ready | (mb_client_tx_err & mb_client_status_we0))) begin
            mb_client_w_pending <= 1'd0;
        end else begin
            mb_client_w_pending <= mb_client_w_pending;
        end
    end
    if (mb_client_status_we0) begin
        mb_client_tx_err <= 1'd0;
    end else begin
        if (((mb_client_wdata_re & (~mb_client_w_ready)) & mb_client_w_pending)) begin
            mb_client_tx_err <= 1'd1;
        end else begin
            mb_client_tx_err <= mb_client_tx_err;
        end
    end
    if (mb_client_status_we0) begin
        mb_client_rx_err <= 1'd0;
    end else begin
        if ((mb_client_rdata_we & (~mb_client_r_valid))) begin
            mb_client_rx_err <= 1'd1;
        end else begin
            mb_client_rx_err <= mb_client_rx_err;
        end
    end
    if (mb_client_available_clear) begin
        mb_client_available_pending <= 1'd0;
    end
    if (mb_client_available_trigger) begin
        mb_client_available_pending <= 1'd1;
    end
    if (mb_client_abort_init_clear) begin
        mb_client_abort_init_pending <= 1'd0;
    end
    mb_client_abort_init_trigger_d <= mb_client_abort_init_trigger;
    if ((mb_client_abort_init_trigger & (~mb_client_abort_init_trigger_d))) begin
        mb_client_abort_init_pending <= 1'd1;
    end
    if (mb_client_abort_done_clear) begin
        mb_client_abort_done_pending <= 1'd0;
    end
    mb_client_abort_done_trigger_d <= mb_client_abort_done_trigger;
    if ((mb_client_abort_done_trigger & (~mb_client_abort_done_trigger_d))) begin
        mb_client_abort_done_pending <= 1'd1;
    end
    if (mb_client_error_clear) begin
        mb_client_error_pending <= 1'd0;
    end
    mb_client_error_trigger_d <= mb_client_error_trigger;
    if ((mb_client_error_trigger & (~mb_client_error_trigger_d))) begin
        mb_client_error_pending <= 1'd1;
    end
    cramsoc_mailboxclient_state <= cramsoc_mailboxclient_next_state;
    if (mb_client_abort_ack1_mailboxclient_next_value_ce0) begin
        mb_client_abort_ack1 <= mb_client_abort_ack1_mailboxclient_next_value0;
    end
    if (mb_client_abort_in_progress1_mailboxclient_next_value_ce1) begin
        mb_client_abort_in_progress1 <= mb_client_abort_in_progress1_mailboxclient_next_value1;
    end
    if (mb_client_w_abort_mailboxclient_next_value_ce2) begin
        mb_client_w_abort <= mb_client_w_abort_mailboxclient_next_value2;
    end
    cramsoc_axilite2csr_state <= cramsoc_axilite2csr_next_state;
    if (cramsoc_last_was_read_axilite2csr_next_value_ce) begin
        cramsoc_last_was_read <= cramsoc_last_was_read_axilite2csr_next_value;
    end
    interface0_bank_bus_dat_r <= 1'd0;
    if (csrbank0_sel) begin
        case (interface0_bank_bus_adr[9:0])
            1'd0: begin
                interface0_bank_bus_dat_r <= csrbank0_control0_w;
            end
            1'd1: begin
                interface0_bank_bus_dat_r <= csrbank0_status_w;
            end
            2'd2: begin
                interface0_bank_bus_dat_r <= csrbank0_map_lo0_w;
            end
            2'd3: begin
                interface0_bank_bus_dat_r <= csrbank0_map_hi0_w;
            end
            3'd4: begin
                interface0_bank_bus_dat_r <= csrbank0_uservalue0_w;
            end
            3'd5: begin
                interface0_bank_bus_dat_r <= csrbank0_protect0_w;
            end
        endcase
    end
    if (csrbank0_control0_re) begin
        coreuser_control_storage[1:0] <= csrbank0_control0_r;
    end
    coreuser_control_re <= csrbank0_control0_re;
    coreuser_status_re <= csrbank0_status_re;
    if (csrbank0_map_lo0_re) begin
        coreuser_map_lo_storage[31:0] <= csrbank0_map_lo0_r;
    end
    coreuser_map_lo_re <= csrbank0_map_lo0_re;
    if (csrbank0_map_hi0_re) begin
        coreuser_map_hi_storage[31:0] <= csrbank0_map_hi0_r;
    end
    coreuser_map_hi_re <= csrbank0_map_hi0_re;
    if (csrbank0_uservalue0_re) begin
        coreuser_uservalue_storage[17:0] <= csrbank0_uservalue0_r;
    end
    coreuser_uservalue_re <= csrbank0_uservalue0_re;
    if (csrbank0_protect0_re) begin
        coreuser_protect_storage <= csrbank0_protect0_r;
    end
    coreuser_protect_re <= csrbank0_protect0_re;
    interface1_bank_bus_dat_r <= 1'd0;
    if (csrbank1_sel) begin
        case (interface1_bank_bus_adr[9:0])
            1'd0: begin
                interface1_bank_bus_dat_r <= csrbank1_wtest0_w;
            end
            1'd1: begin
                interface1_bank_bus_dat_r <= csrbank1_rtest_w;
            end
        endcase
    end
    if (csrbank1_wtest0_re) begin
        csr_wtest_storage[31:0] <= csrbank1_wtest0_r;
    end
    csr_wtest_re <= csrbank1_wtest0_re;
    csr_rtest_re <= csrbank1_rtest_re;
    interface2_bank_bus_dat_r <= 1'd0;
    if (csrbank2_sel) begin
        case (interface2_bank_bus_adr[9:0])
            1'd0: begin
                interface2_bank_bus_dat_r <= csrbank2_control0_w;
            end
            1'd1: begin
                interface2_bank_bus_dat_r <= csrbank2_heartbeat_w;
            end
        endcase
    end
    if (csrbank2_control0_re) begin
        d11ctime_control_storage[31:0] <= csrbank2_control0_r;
    end
    d11ctime_control_re <= csrbank2_control0_re;
    d11ctime_heartbeat_re <= csrbank2_heartbeat_re;
    interface3_bank_bus_dat_r <= 1'd0;
    if (csrbank3_sel) begin
        case (interface3_bank_bus_adr[9:0])
            1'd0: begin
                interface3_bank_bus_dat_r <= csrbank3_ev_soft0_w;
            end
            1'd1: begin
                interface3_bank_bus_dat_r <= csrbank3_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface3_bank_bus_dat_r <= csrbank3_ev_polarity0_w;
            end
            2'd3: begin
                interface3_bank_bus_dat_r <= csrbank3_ev_status_w;
            end
            3'd4: begin
                interface3_bank_bus_dat_r <= csrbank3_ev_pending_w;
            end
            3'd5: begin
                interface3_bank_bus_dat_r <= csrbank3_ev_enable0_w;
            end
        endcase
    end
    if (csrbank3_ev_soft0_re) begin
        irqarray0_soft_storage[15:0] <= csrbank3_ev_soft0_r;
    end
    irqarray0_soft_re <= csrbank3_ev_soft0_re;
    if (csrbank3_ev_edge_triggered0_re) begin
        irqarray0_edge_triggered_storage[15:0] <= csrbank3_ev_edge_triggered0_r;
    end
    irqarray0_edge_triggered_re <= csrbank3_ev_edge_triggered0_re;
    if (csrbank3_ev_polarity0_re) begin
        irqarray0_polarity_storage[15:0] <= csrbank3_ev_polarity0_r;
    end
    irqarray0_polarity_re <= csrbank3_ev_polarity0_re;
    irqarray0_status_re <= csrbank3_ev_status_re;
    if (csrbank3_ev_pending_re) begin
        irqarray0_pending_r[15:0] <= csrbank3_ev_pending_r;
    end
    irqarray0_pending_re <= csrbank3_ev_pending_re;
    if (csrbank3_ev_enable0_re) begin
        irqarray0_enable_storage[15:0] <= csrbank3_ev_enable0_r;
    end
    irqarray0_enable_re <= csrbank3_ev_enable0_re;
    interface4_bank_bus_dat_r <= 1'd0;
    if (csrbank4_sel) begin
        case (interface4_bank_bus_adr[9:0])
            1'd0: begin
                interface4_bank_bus_dat_r <= csrbank4_ev_soft0_w;
            end
            1'd1: begin
                interface4_bank_bus_dat_r <= csrbank4_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface4_bank_bus_dat_r <= csrbank4_ev_polarity0_w;
            end
            2'd3: begin
                interface4_bank_bus_dat_r <= csrbank4_ev_status_w;
            end
            3'd4: begin
                interface4_bank_bus_dat_r <= csrbank4_ev_pending_w;
            end
            3'd5: begin
                interface4_bank_bus_dat_r <= csrbank4_ev_enable0_w;
            end
        endcase
    end
    if (csrbank4_ev_soft0_re) begin
        irqarray1_soft_storage[15:0] <= csrbank4_ev_soft0_r;
    end
    irqarray1_soft_re <= csrbank4_ev_soft0_re;
    if (csrbank4_ev_edge_triggered0_re) begin
        irqarray1_edge_triggered_storage[15:0] <= csrbank4_ev_edge_triggered0_r;
    end
    irqarray1_edge_triggered_re <= csrbank4_ev_edge_triggered0_re;
    if (csrbank4_ev_polarity0_re) begin
        irqarray1_polarity_storage[15:0] <= csrbank4_ev_polarity0_r;
    end
    irqarray1_polarity_re <= csrbank4_ev_polarity0_re;
    irqarray1_status_re <= csrbank4_ev_status_re;
    if (csrbank4_ev_pending_re) begin
        irqarray1_pending_r[15:0] <= csrbank4_ev_pending_r;
    end
    irqarray1_pending_re <= csrbank4_ev_pending_re;
    if (csrbank4_ev_enable0_re) begin
        irqarray1_enable_storage[15:0] <= csrbank4_ev_enable0_r;
    end
    irqarray1_enable_re <= csrbank4_ev_enable0_re;
    interface5_bank_bus_dat_r <= 1'd0;
    if (csrbank5_sel) begin
        case (interface5_bank_bus_adr[9:0])
            1'd0: begin
                interface5_bank_bus_dat_r <= csrbank5_ev_soft0_w;
            end
            1'd1: begin
                interface5_bank_bus_dat_r <= csrbank5_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface5_bank_bus_dat_r <= csrbank5_ev_polarity0_w;
            end
            2'd3: begin
                interface5_bank_bus_dat_r <= csrbank5_ev_status_w;
            end
            3'd4: begin
                interface5_bank_bus_dat_r <= csrbank5_ev_pending_w;
            end
            3'd5: begin
                interface5_bank_bus_dat_r <= csrbank5_ev_enable0_w;
            end
        endcase
    end
    if (csrbank5_ev_soft0_re) begin
        irqarray10_soft_storage[15:0] <= csrbank5_ev_soft0_r;
    end
    irqarray10_soft_re <= csrbank5_ev_soft0_re;
    if (csrbank5_ev_edge_triggered0_re) begin
        irqarray10_edge_triggered_storage[15:0] <= csrbank5_ev_edge_triggered0_r;
    end
    irqarray10_edge_triggered_re <= csrbank5_ev_edge_triggered0_re;
    if (csrbank5_ev_polarity0_re) begin
        irqarray10_polarity_storage[15:0] <= csrbank5_ev_polarity0_r;
    end
    irqarray10_polarity_re <= csrbank5_ev_polarity0_re;
    irqarray10_status_re <= csrbank5_ev_status_re;
    if (csrbank5_ev_pending_re) begin
        irqarray10_pending_r[15:0] <= csrbank5_ev_pending_r;
    end
    irqarray10_pending_re <= csrbank5_ev_pending_re;
    if (csrbank5_ev_enable0_re) begin
        irqarray10_enable_storage[15:0] <= csrbank5_ev_enable0_r;
    end
    irqarray10_enable_re <= csrbank5_ev_enable0_re;
    interface6_bank_bus_dat_r <= 1'd0;
    if (csrbank6_sel) begin
        case (interface6_bank_bus_adr[9:0])
            1'd0: begin
                interface6_bank_bus_dat_r <= csrbank6_ev_soft0_w;
            end
            1'd1: begin
                interface6_bank_bus_dat_r <= csrbank6_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface6_bank_bus_dat_r <= csrbank6_ev_polarity0_w;
            end
            2'd3: begin
                interface6_bank_bus_dat_r <= csrbank6_ev_status_w;
            end
            3'd4: begin
                interface6_bank_bus_dat_r <= csrbank6_ev_pending_w;
            end
            3'd5: begin
                interface6_bank_bus_dat_r <= csrbank6_ev_enable0_w;
            end
        endcase
    end
    if (csrbank6_ev_soft0_re) begin
        irqarray11_soft_storage[15:0] <= csrbank6_ev_soft0_r;
    end
    irqarray11_soft_re <= csrbank6_ev_soft0_re;
    if (csrbank6_ev_edge_triggered0_re) begin
        irqarray11_edge_triggered_storage[15:0] <= csrbank6_ev_edge_triggered0_r;
    end
    irqarray11_edge_triggered_re <= csrbank6_ev_edge_triggered0_re;
    if (csrbank6_ev_polarity0_re) begin
        irqarray11_polarity_storage[15:0] <= csrbank6_ev_polarity0_r;
    end
    irqarray11_polarity_re <= csrbank6_ev_polarity0_re;
    irqarray11_status_re <= csrbank6_ev_status_re;
    if (csrbank6_ev_pending_re) begin
        irqarray11_pending_r[15:0] <= csrbank6_ev_pending_r;
    end
    irqarray11_pending_re <= csrbank6_ev_pending_re;
    if (csrbank6_ev_enable0_re) begin
        irqarray11_enable_storage[15:0] <= csrbank6_ev_enable0_r;
    end
    irqarray11_enable_re <= csrbank6_ev_enable0_re;
    interface7_bank_bus_dat_r <= 1'd0;
    if (csrbank7_sel) begin
        case (interface7_bank_bus_adr[9:0])
            1'd0: begin
                interface7_bank_bus_dat_r <= csrbank7_ev_soft0_w;
            end
            1'd1: begin
                interface7_bank_bus_dat_r <= csrbank7_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface7_bank_bus_dat_r <= csrbank7_ev_polarity0_w;
            end
            2'd3: begin
                interface7_bank_bus_dat_r <= csrbank7_ev_status_w;
            end
            3'd4: begin
                interface7_bank_bus_dat_r <= csrbank7_ev_pending_w;
            end
            3'd5: begin
                interface7_bank_bus_dat_r <= csrbank7_ev_enable0_w;
            end
        endcase
    end
    if (csrbank7_ev_soft0_re) begin
        irqarray12_soft_storage[15:0] <= csrbank7_ev_soft0_r;
    end
    irqarray12_soft_re <= csrbank7_ev_soft0_re;
    if (csrbank7_ev_edge_triggered0_re) begin
        irqarray12_edge_triggered_storage[15:0] <= csrbank7_ev_edge_triggered0_r;
    end
    irqarray12_edge_triggered_re <= csrbank7_ev_edge_triggered0_re;
    if (csrbank7_ev_polarity0_re) begin
        irqarray12_polarity_storage[15:0] <= csrbank7_ev_polarity0_r;
    end
    irqarray12_polarity_re <= csrbank7_ev_polarity0_re;
    irqarray12_status_re <= csrbank7_ev_status_re;
    if (csrbank7_ev_pending_re) begin
        irqarray12_pending_r[15:0] <= csrbank7_ev_pending_r;
    end
    irqarray12_pending_re <= csrbank7_ev_pending_re;
    if (csrbank7_ev_enable0_re) begin
        irqarray12_enable_storage[15:0] <= csrbank7_ev_enable0_r;
    end
    irqarray12_enable_re <= csrbank7_ev_enable0_re;
    interface8_bank_bus_dat_r <= 1'd0;
    if (csrbank8_sel) begin
        case (interface8_bank_bus_adr[9:0])
            1'd0: begin
                interface8_bank_bus_dat_r <= csrbank8_ev_soft0_w;
            end
            1'd1: begin
                interface8_bank_bus_dat_r <= csrbank8_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface8_bank_bus_dat_r <= csrbank8_ev_polarity0_w;
            end
            2'd3: begin
                interface8_bank_bus_dat_r <= csrbank8_ev_status_w;
            end
            3'd4: begin
                interface8_bank_bus_dat_r <= csrbank8_ev_pending_w;
            end
            3'd5: begin
                interface8_bank_bus_dat_r <= csrbank8_ev_enable0_w;
            end
        endcase
    end
    if (csrbank8_ev_soft0_re) begin
        irqarray13_soft_storage[15:0] <= csrbank8_ev_soft0_r;
    end
    irqarray13_soft_re <= csrbank8_ev_soft0_re;
    if (csrbank8_ev_edge_triggered0_re) begin
        irqarray13_edge_triggered_storage[15:0] <= csrbank8_ev_edge_triggered0_r;
    end
    irqarray13_edge_triggered_re <= csrbank8_ev_edge_triggered0_re;
    if (csrbank8_ev_polarity0_re) begin
        irqarray13_polarity_storage[15:0] <= csrbank8_ev_polarity0_r;
    end
    irqarray13_polarity_re <= csrbank8_ev_polarity0_re;
    irqarray13_status_re <= csrbank8_ev_status_re;
    if (csrbank8_ev_pending_re) begin
        irqarray13_pending_r[15:0] <= csrbank8_ev_pending_r;
    end
    irqarray13_pending_re <= csrbank8_ev_pending_re;
    if (csrbank8_ev_enable0_re) begin
        irqarray13_enable_storage[15:0] <= csrbank8_ev_enable0_r;
    end
    irqarray13_enable_re <= csrbank8_ev_enable0_re;
    interface9_bank_bus_dat_r <= 1'd0;
    if (csrbank9_sel) begin
        case (interface9_bank_bus_adr[9:0])
            1'd0: begin
                interface9_bank_bus_dat_r <= csrbank9_ev_soft0_w;
            end
            1'd1: begin
                interface9_bank_bus_dat_r <= csrbank9_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface9_bank_bus_dat_r <= csrbank9_ev_polarity0_w;
            end
            2'd3: begin
                interface9_bank_bus_dat_r <= csrbank9_ev_status_w;
            end
            3'd4: begin
                interface9_bank_bus_dat_r <= csrbank9_ev_pending_w;
            end
            3'd5: begin
                interface9_bank_bus_dat_r <= csrbank9_ev_enable0_w;
            end
        endcase
    end
    if (csrbank9_ev_soft0_re) begin
        irqarray14_soft_storage[15:0] <= csrbank9_ev_soft0_r;
    end
    irqarray14_soft_re <= csrbank9_ev_soft0_re;
    if (csrbank9_ev_edge_triggered0_re) begin
        irqarray14_edge_triggered_storage[15:0] <= csrbank9_ev_edge_triggered0_r;
    end
    irqarray14_edge_triggered_re <= csrbank9_ev_edge_triggered0_re;
    if (csrbank9_ev_polarity0_re) begin
        irqarray14_polarity_storage[15:0] <= csrbank9_ev_polarity0_r;
    end
    irqarray14_polarity_re <= csrbank9_ev_polarity0_re;
    irqarray14_status_re <= csrbank9_ev_status_re;
    if (csrbank9_ev_pending_re) begin
        irqarray14_pending_r[15:0] <= csrbank9_ev_pending_r;
    end
    irqarray14_pending_re <= csrbank9_ev_pending_re;
    if (csrbank9_ev_enable0_re) begin
        irqarray14_enable_storage[15:0] <= csrbank9_ev_enable0_r;
    end
    irqarray14_enable_re <= csrbank9_ev_enable0_re;
    interface10_bank_bus_dat_r <= 1'd0;
    if (csrbank10_sel) begin
        case (interface10_bank_bus_adr[9:0])
            1'd0: begin
                interface10_bank_bus_dat_r <= csrbank10_ev_soft0_w;
            end
            1'd1: begin
                interface10_bank_bus_dat_r <= csrbank10_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface10_bank_bus_dat_r <= csrbank10_ev_polarity0_w;
            end
            2'd3: begin
                interface10_bank_bus_dat_r <= csrbank10_ev_status_w;
            end
            3'd4: begin
                interface10_bank_bus_dat_r <= csrbank10_ev_pending_w;
            end
            3'd5: begin
                interface10_bank_bus_dat_r <= csrbank10_ev_enable0_w;
            end
        endcase
    end
    if (csrbank10_ev_soft0_re) begin
        irqarray15_soft_storage[15:0] <= csrbank10_ev_soft0_r;
    end
    irqarray15_soft_re <= csrbank10_ev_soft0_re;
    if (csrbank10_ev_edge_triggered0_re) begin
        irqarray15_edge_triggered_storage[15:0] <= csrbank10_ev_edge_triggered0_r;
    end
    irqarray15_edge_triggered_re <= csrbank10_ev_edge_triggered0_re;
    if (csrbank10_ev_polarity0_re) begin
        irqarray15_polarity_storage[15:0] <= csrbank10_ev_polarity0_r;
    end
    irqarray15_polarity_re <= csrbank10_ev_polarity0_re;
    irqarray15_status_re <= csrbank10_ev_status_re;
    if (csrbank10_ev_pending_re) begin
        irqarray15_pending_r[15:0] <= csrbank10_ev_pending_r;
    end
    irqarray15_pending_re <= csrbank10_ev_pending_re;
    if (csrbank10_ev_enable0_re) begin
        irqarray15_enable_storage[15:0] <= csrbank10_ev_enable0_r;
    end
    irqarray15_enable_re <= csrbank10_ev_enable0_re;
    interface11_bank_bus_dat_r <= 1'd0;
    if (csrbank11_sel) begin
        case (interface11_bank_bus_adr[9:0])
            1'd0: begin
                interface11_bank_bus_dat_r <= csrbank11_ev_soft0_w;
            end
            1'd1: begin
                interface11_bank_bus_dat_r <= csrbank11_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface11_bank_bus_dat_r <= csrbank11_ev_polarity0_w;
            end
            2'd3: begin
                interface11_bank_bus_dat_r <= csrbank11_ev_status_w;
            end
            3'd4: begin
                interface11_bank_bus_dat_r <= csrbank11_ev_pending_w;
            end
            3'd5: begin
                interface11_bank_bus_dat_r <= csrbank11_ev_enable0_w;
            end
        endcase
    end
    if (csrbank11_ev_soft0_re) begin
        irqarray16_soft_storage[15:0] <= csrbank11_ev_soft0_r;
    end
    irqarray16_soft_re <= csrbank11_ev_soft0_re;
    if (csrbank11_ev_edge_triggered0_re) begin
        irqarray16_edge_triggered_storage[15:0] <= csrbank11_ev_edge_triggered0_r;
    end
    irqarray16_edge_triggered_re <= csrbank11_ev_edge_triggered0_re;
    if (csrbank11_ev_polarity0_re) begin
        irqarray16_polarity_storage[15:0] <= csrbank11_ev_polarity0_r;
    end
    irqarray16_polarity_re <= csrbank11_ev_polarity0_re;
    irqarray16_status_re <= csrbank11_ev_status_re;
    if (csrbank11_ev_pending_re) begin
        irqarray16_pending_r[15:0] <= csrbank11_ev_pending_r;
    end
    irqarray16_pending_re <= csrbank11_ev_pending_re;
    if (csrbank11_ev_enable0_re) begin
        irqarray16_enable_storage[15:0] <= csrbank11_ev_enable0_r;
    end
    irqarray16_enable_re <= csrbank11_ev_enable0_re;
    interface12_bank_bus_dat_r <= 1'd0;
    if (csrbank12_sel) begin
        case (interface12_bank_bus_adr[9:0])
            1'd0: begin
                interface12_bank_bus_dat_r <= csrbank12_ev_soft0_w;
            end
            1'd1: begin
                interface12_bank_bus_dat_r <= csrbank12_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface12_bank_bus_dat_r <= csrbank12_ev_polarity0_w;
            end
            2'd3: begin
                interface12_bank_bus_dat_r <= csrbank12_ev_status_w;
            end
            3'd4: begin
                interface12_bank_bus_dat_r <= csrbank12_ev_pending_w;
            end
            3'd5: begin
                interface12_bank_bus_dat_r <= csrbank12_ev_enable0_w;
            end
        endcase
    end
    if (csrbank12_ev_soft0_re) begin
        irqarray17_soft_storage[15:0] <= csrbank12_ev_soft0_r;
    end
    irqarray17_soft_re <= csrbank12_ev_soft0_re;
    if (csrbank12_ev_edge_triggered0_re) begin
        irqarray17_edge_triggered_storage[15:0] <= csrbank12_ev_edge_triggered0_r;
    end
    irqarray17_edge_triggered_re <= csrbank12_ev_edge_triggered0_re;
    if (csrbank12_ev_polarity0_re) begin
        irqarray17_polarity_storage[15:0] <= csrbank12_ev_polarity0_r;
    end
    irqarray17_polarity_re <= csrbank12_ev_polarity0_re;
    irqarray17_status_re <= csrbank12_ev_status_re;
    if (csrbank12_ev_pending_re) begin
        irqarray17_pending_r[15:0] <= csrbank12_ev_pending_r;
    end
    irqarray17_pending_re <= csrbank12_ev_pending_re;
    if (csrbank12_ev_enable0_re) begin
        irqarray17_enable_storage[15:0] <= csrbank12_ev_enable0_r;
    end
    irqarray17_enable_re <= csrbank12_ev_enable0_re;
    interface13_bank_bus_dat_r <= 1'd0;
    if (csrbank13_sel) begin
        case (interface13_bank_bus_adr[9:0])
            1'd0: begin
                interface13_bank_bus_dat_r <= csrbank13_ev_soft0_w;
            end
            1'd1: begin
                interface13_bank_bus_dat_r <= csrbank13_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface13_bank_bus_dat_r <= csrbank13_ev_polarity0_w;
            end
            2'd3: begin
                interface13_bank_bus_dat_r <= csrbank13_ev_status_w;
            end
            3'd4: begin
                interface13_bank_bus_dat_r <= csrbank13_ev_pending_w;
            end
            3'd5: begin
                interface13_bank_bus_dat_r <= csrbank13_ev_enable0_w;
            end
        endcase
    end
    if (csrbank13_ev_soft0_re) begin
        irqarray18_soft_storage[15:0] <= csrbank13_ev_soft0_r;
    end
    irqarray18_soft_re <= csrbank13_ev_soft0_re;
    if (csrbank13_ev_edge_triggered0_re) begin
        irqarray18_edge_triggered_storage[15:0] <= csrbank13_ev_edge_triggered0_r;
    end
    irqarray18_edge_triggered_re <= csrbank13_ev_edge_triggered0_re;
    if (csrbank13_ev_polarity0_re) begin
        irqarray18_polarity_storage[15:0] <= csrbank13_ev_polarity0_r;
    end
    irqarray18_polarity_re <= csrbank13_ev_polarity0_re;
    irqarray18_status_re <= csrbank13_ev_status_re;
    if (csrbank13_ev_pending_re) begin
        irqarray18_pending_r[15:0] <= csrbank13_ev_pending_r;
    end
    irqarray18_pending_re <= csrbank13_ev_pending_re;
    if (csrbank13_ev_enable0_re) begin
        irqarray18_enable_storage[15:0] <= csrbank13_ev_enable0_r;
    end
    irqarray18_enable_re <= csrbank13_ev_enable0_re;
    interface14_bank_bus_dat_r <= 1'd0;
    if (csrbank14_sel) begin
        case (interface14_bank_bus_adr[9:0])
            1'd0: begin
                interface14_bank_bus_dat_r <= csrbank14_ev_soft0_w;
            end
            1'd1: begin
                interface14_bank_bus_dat_r <= csrbank14_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface14_bank_bus_dat_r <= csrbank14_ev_polarity0_w;
            end
            2'd3: begin
                interface14_bank_bus_dat_r <= csrbank14_ev_status_w;
            end
            3'd4: begin
                interface14_bank_bus_dat_r <= csrbank14_ev_pending_w;
            end
            3'd5: begin
                interface14_bank_bus_dat_r <= csrbank14_ev_enable0_w;
            end
        endcase
    end
    if (csrbank14_ev_soft0_re) begin
        irqarray19_soft_storage[15:0] <= csrbank14_ev_soft0_r;
    end
    irqarray19_soft_re <= csrbank14_ev_soft0_re;
    if (csrbank14_ev_edge_triggered0_re) begin
        irqarray19_edge_triggered_storage[15:0] <= csrbank14_ev_edge_triggered0_r;
    end
    irqarray19_edge_triggered_re <= csrbank14_ev_edge_triggered0_re;
    if (csrbank14_ev_polarity0_re) begin
        irqarray19_polarity_storage[15:0] <= csrbank14_ev_polarity0_r;
    end
    irqarray19_polarity_re <= csrbank14_ev_polarity0_re;
    irqarray19_status_re <= csrbank14_ev_status_re;
    if (csrbank14_ev_pending_re) begin
        irqarray19_pending_r[15:0] <= csrbank14_ev_pending_r;
    end
    irqarray19_pending_re <= csrbank14_ev_pending_re;
    if (csrbank14_ev_enable0_re) begin
        irqarray19_enable_storage[15:0] <= csrbank14_ev_enable0_r;
    end
    irqarray19_enable_re <= csrbank14_ev_enable0_re;
    interface15_bank_bus_dat_r <= 1'd0;
    if (csrbank15_sel) begin
        case (interface15_bank_bus_adr[9:0])
            1'd0: begin
                interface15_bank_bus_dat_r <= csrbank15_ev_soft0_w;
            end
            1'd1: begin
                interface15_bank_bus_dat_r <= csrbank15_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface15_bank_bus_dat_r <= csrbank15_ev_polarity0_w;
            end
            2'd3: begin
                interface15_bank_bus_dat_r <= csrbank15_ev_status_w;
            end
            3'd4: begin
                interface15_bank_bus_dat_r <= csrbank15_ev_pending_w;
            end
            3'd5: begin
                interface15_bank_bus_dat_r <= csrbank15_ev_enable0_w;
            end
        endcase
    end
    if (csrbank15_ev_soft0_re) begin
        irqarray2_soft_storage[15:0] <= csrbank15_ev_soft0_r;
    end
    irqarray2_soft_re <= csrbank15_ev_soft0_re;
    if (csrbank15_ev_edge_triggered0_re) begin
        irqarray2_edge_triggered_storage[15:0] <= csrbank15_ev_edge_triggered0_r;
    end
    irqarray2_edge_triggered_re <= csrbank15_ev_edge_triggered0_re;
    if (csrbank15_ev_polarity0_re) begin
        irqarray2_polarity_storage[15:0] <= csrbank15_ev_polarity0_r;
    end
    irqarray2_polarity_re <= csrbank15_ev_polarity0_re;
    irqarray2_status_re <= csrbank15_ev_status_re;
    if (csrbank15_ev_pending_re) begin
        irqarray2_pending_r[15:0] <= csrbank15_ev_pending_r;
    end
    irqarray2_pending_re <= csrbank15_ev_pending_re;
    if (csrbank15_ev_enable0_re) begin
        irqarray2_enable_storage[15:0] <= csrbank15_ev_enable0_r;
    end
    irqarray2_enable_re <= csrbank15_ev_enable0_re;
    interface16_bank_bus_dat_r <= 1'd0;
    if (csrbank16_sel) begin
        case (interface16_bank_bus_adr[9:0])
            1'd0: begin
                interface16_bank_bus_dat_r <= csrbank16_ev_soft0_w;
            end
            1'd1: begin
                interface16_bank_bus_dat_r <= csrbank16_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface16_bank_bus_dat_r <= csrbank16_ev_polarity0_w;
            end
            2'd3: begin
                interface16_bank_bus_dat_r <= csrbank16_ev_status_w;
            end
            3'd4: begin
                interface16_bank_bus_dat_r <= csrbank16_ev_pending_w;
            end
            3'd5: begin
                interface16_bank_bus_dat_r <= csrbank16_ev_enable0_w;
            end
        endcase
    end
    if (csrbank16_ev_soft0_re) begin
        irqarray3_soft_storage[15:0] <= csrbank16_ev_soft0_r;
    end
    irqarray3_soft_re <= csrbank16_ev_soft0_re;
    if (csrbank16_ev_edge_triggered0_re) begin
        irqarray3_edge_triggered_storage[15:0] <= csrbank16_ev_edge_triggered0_r;
    end
    irqarray3_edge_triggered_re <= csrbank16_ev_edge_triggered0_re;
    if (csrbank16_ev_polarity0_re) begin
        irqarray3_polarity_storage[15:0] <= csrbank16_ev_polarity0_r;
    end
    irqarray3_polarity_re <= csrbank16_ev_polarity0_re;
    irqarray3_status_re <= csrbank16_ev_status_re;
    if (csrbank16_ev_pending_re) begin
        irqarray3_pending_r[15:0] <= csrbank16_ev_pending_r;
    end
    irqarray3_pending_re <= csrbank16_ev_pending_re;
    if (csrbank16_ev_enable0_re) begin
        irqarray3_enable_storage[15:0] <= csrbank16_ev_enable0_r;
    end
    irqarray3_enable_re <= csrbank16_ev_enable0_re;
    interface17_bank_bus_dat_r <= 1'd0;
    if (csrbank17_sel) begin
        case (interface17_bank_bus_adr[9:0])
            1'd0: begin
                interface17_bank_bus_dat_r <= csrbank17_ev_soft0_w;
            end
            1'd1: begin
                interface17_bank_bus_dat_r <= csrbank17_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface17_bank_bus_dat_r <= csrbank17_ev_polarity0_w;
            end
            2'd3: begin
                interface17_bank_bus_dat_r <= csrbank17_ev_status_w;
            end
            3'd4: begin
                interface17_bank_bus_dat_r <= csrbank17_ev_pending_w;
            end
            3'd5: begin
                interface17_bank_bus_dat_r <= csrbank17_ev_enable0_w;
            end
        endcase
    end
    if (csrbank17_ev_soft0_re) begin
        irqarray4_soft_storage[15:0] <= csrbank17_ev_soft0_r;
    end
    irqarray4_soft_re <= csrbank17_ev_soft0_re;
    if (csrbank17_ev_edge_triggered0_re) begin
        irqarray4_edge_triggered_storage[15:0] <= csrbank17_ev_edge_triggered0_r;
    end
    irqarray4_edge_triggered_re <= csrbank17_ev_edge_triggered0_re;
    if (csrbank17_ev_polarity0_re) begin
        irqarray4_polarity_storage[15:0] <= csrbank17_ev_polarity0_r;
    end
    irqarray4_polarity_re <= csrbank17_ev_polarity0_re;
    irqarray4_status_re <= csrbank17_ev_status_re;
    if (csrbank17_ev_pending_re) begin
        irqarray4_pending_r[15:0] <= csrbank17_ev_pending_r;
    end
    irqarray4_pending_re <= csrbank17_ev_pending_re;
    if (csrbank17_ev_enable0_re) begin
        irqarray4_enable_storage[15:0] <= csrbank17_ev_enable0_r;
    end
    irqarray4_enable_re <= csrbank17_ev_enable0_re;
    interface18_bank_bus_dat_r <= 1'd0;
    if (csrbank18_sel) begin
        case (interface18_bank_bus_adr[9:0])
            1'd0: begin
                interface18_bank_bus_dat_r <= csrbank18_ev_soft0_w;
            end
            1'd1: begin
                interface18_bank_bus_dat_r <= csrbank18_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface18_bank_bus_dat_r <= csrbank18_ev_polarity0_w;
            end
            2'd3: begin
                interface18_bank_bus_dat_r <= csrbank18_ev_status_w;
            end
            3'd4: begin
                interface18_bank_bus_dat_r <= csrbank18_ev_pending_w;
            end
            3'd5: begin
                interface18_bank_bus_dat_r <= csrbank18_ev_enable0_w;
            end
        endcase
    end
    if (csrbank18_ev_soft0_re) begin
        irqarray5_soft_storage[15:0] <= csrbank18_ev_soft0_r;
    end
    irqarray5_soft_re <= csrbank18_ev_soft0_re;
    if (csrbank18_ev_edge_triggered0_re) begin
        irqarray5_edge_triggered_storage[15:0] <= csrbank18_ev_edge_triggered0_r;
    end
    irqarray5_edge_triggered_re <= csrbank18_ev_edge_triggered0_re;
    if (csrbank18_ev_polarity0_re) begin
        irqarray5_polarity_storage[15:0] <= csrbank18_ev_polarity0_r;
    end
    irqarray5_polarity_re <= csrbank18_ev_polarity0_re;
    irqarray5_status_re <= csrbank18_ev_status_re;
    if (csrbank18_ev_pending_re) begin
        irqarray5_pending_r[15:0] <= csrbank18_ev_pending_r;
    end
    irqarray5_pending_re <= csrbank18_ev_pending_re;
    if (csrbank18_ev_enable0_re) begin
        irqarray5_enable_storage[15:0] <= csrbank18_ev_enable0_r;
    end
    irqarray5_enable_re <= csrbank18_ev_enable0_re;
    interface19_bank_bus_dat_r <= 1'd0;
    if (csrbank19_sel) begin
        case (interface19_bank_bus_adr[9:0])
            1'd0: begin
                interface19_bank_bus_dat_r <= csrbank19_ev_soft0_w;
            end
            1'd1: begin
                interface19_bank_bus_dat_r <= csrbank19_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface19_bank_bus_dat_r <= csrbank19_ev_polarity0_w;
            end
            2'd3: begin
                interface19_bank_bus_dat_r <= csrbank19_ev_status_w;
            end
            3'd4: begin
                interface19_bank_bus_dat_r <= csrbank19_ev_pending_w;
            end
            3'd5: begin
                interface19_bank_bus_dat_r <= csrbank19_ev_enable0_w;
            end
        endcase
    end
    if (csrbank19_ev_soft0_re) begin
        irqarray6_soft_storage[15:0] <= csrbank19_ev_soft0_r;
    end
    irqarray6_soft_re <= csrbank19_ev_soft0_re;
    if (csrbank19_ev_edge_triggered0_re) begin
        irqarray6_edge_triggered_storage[15:0] <= csrbank19_ev_edge_triggered0_r;
    end
    irqarray6_edge_triggered_re <= csrbank19_ev_edge_triggered0_re;
    if (csrbank19_ev_polarity0_re) begin
        irqarray6_polarity_storage[15:0] <= csrbank19_ev_polarity0_r;
    end
    irqarray6_polarity_re <= csrbank19_ev_polarity0_re;
    irqarray6_status_re <= csrbank19_ev_status_re;
    if (csrbank19_ev_pending_re) begin
        irqarray6_pending_r[15:0] <= csrbank19_ev_pending_r;
    end
    irqarray6_pending_re <= csrbank19_ev_pending_re;
    if (csrbank19_ev_enable0_re) begin
        irqarray6_enable_storage[15:0] <= csrbank19_ev_enable0_r;
    end
    irqarray6_enable_re <= csrbank19_ev_enable0_re;
    interface20_bank_bus_dat_r <= 1'd0;
    if (csrbank20_sel) begin
        case (interface20_bank_bus_adr[9:0])
            1'd0: begin
                interface20_bank_bus_dat_r <= csrbank20_ev_soft0_w;
            end
            1'd1: begin
                interface20_bank_bus_dat_r <= csrbank20_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface20_bank_bus_dat_r <= csrbank20_ev_polarity0_w;
            end
            2'd3: begin
                interface20_bank_bus_dat_r <= csrbank20_ev_status_w;
            end
            3'd4: begin
                interface20_bank_bus_dat_r <= csrbank20_ev_pending_w;
            end
            3'd5: begin
                interface20_bank_bus_dat_r <= csrbank20_ev_enable0_w;
            end
        endcase
    end
    if (csrbank20_ev_soft0_re) begin
        irqarray7_soft_storage[15:0] <= csrbank20_ev_soft0_r;
    end
    irqarray7_soft_re <= csrbank20_ev_soft0_re;
    if (csrbank20_ev_edge_triggered0_re) begin
        irqarray7_edge_triggered_storage[15:0] <= csrbank20_ev_edge_triggered0_r;
    end
    irqarray7_edge_triggered_re <= csrbank20_ev_edge_triggered0_re;
    if (csrbank20_ev_polarity0_re) begin
        irqarray7_polarity_storage[15:0] <= csrbank20_ev_polarity0_r;
    end
    irqarray7_polarity_re <= csrbank20_ev_polarity0_re;
    irqarray7_status_re <= csrbank20_ev_status_re;
    if (csrbank20_ev_pending_re) begin
        irqarray7_pending_r[15:0] <= csrbank20_ev_pending_r;
    end
    irqarray7_pending_re <= csrbank20_ev_pending_re;
    if (csrbank20_ev_enable0_re) begin
        irqarray7_enable_storage[15:0] <= csrbank20_ev_enable0_r;
    end
    irqarray7_enable_re <= csrbank20_ev_enable0_re;
    interface21_bank_bus_dat_r <= 1'd0;
    if (csrbank21_sel) begin
        case (interface21_bank_bus_adr[9:0])
            1'd0: begin
                interface21_bank_bus_dat_r <= csrbank21_ev_soft0_w;
            end
            1'd1: begin
                interface21_bank_bus_dat_r <= csrbank21_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface21_bank_bus_dat_r <= csrbank21_ev_polarity0_w;
            end
            2'd3: begin
                interface21_bank_bus_dat_r <= csrbank21_ev_status_w;
            end
            3'd4: begin
                interface21_bank_bus_dat_r <= csrbank21_ev_pending_w;
            end
            3'd5: begin
                interface21_bank_bus_dat_r <= csrbank21_ev_enable0_w;
            end
        endcase
    end
    if (csrbank21_ev_soft0_re) begin
        irqarray8_soft_storage[15:0] <= csrbank21_ev_soft0_r;
    end
    irqarray8_soft_re <= csrbank21_ev_soft0_re;
    if (csrbank21_ev_edge_triggered0_re) begin
        irqarray8_edge_triggered_storage[15:0] <= csrbank21_ev_edge_triggered0_r;
    end
    irqarray8_edge_triggered_re <= csrbank21_ev_edge_triggered0_re;
    if (csrbank21_ev_polarity0_re) begin
        irqarray8_polarity_storage[15:0] <= csrbank21_ev_polarity0_r;
    end
    irqarray8_polarity_re <= csrbank21_ev_polarity0_re;
    irqarray8_status_re <= csrbank21_ev_status_re;
    if (csrbank21_ev_pending_re) begin
        irqarray8_pending_r[15:0] <= csrbank21_ev_pending_r;
    end
    irqarray8_pending_re <= csrbank21_ev_pending_re;
    if (csrbank21_ev_enable0_re) begin
        irqarray8_enable_storage[15:0] <= csrbank21_ev_enable0_r;
    end
    irqarray8_enable_re <= csrbank21_ev_enable0_re;
    interface22_bank_bus_dat_r <= 1'd0;
    if (csrbank22_sel) begin
        case (interface22_bank_bus_adr[9:0])
            1'd0: begin
                interface22_bank_bus_dat_r <= csrbank22_ev_soft0_w;
            end
            1'd1: begin
                interface22_bank_bus_dat_r <= csrbank22_ev_edge_triggered0_w;
            end
            2'd2: begin
                interface22_bank_bus_dat_r <= csrbank22_ev_polarity0_w;
            end
            2'd3: begin
                interface22_bank_bus_dat_r <= csrbank22_ev_status_w;
            end
            3'd4: begin
                interface22_bank_bus_dat_r <= csrbank22_ev_pending_w;
            end
            3'd5: begin
                interface22_bank_bus_dat_r <= csrbank22_ev_enable0_w;
            end
        endcase
    end
    if (csrbank22_ev_soft0_re) begin
        irqarray9_soft_storage[15:0] <= csrbank22_ev_soft0_r;
    end
    irqarray9_soft_re <= csrbank22_ev_soft0_re;
    if (csrbank22_ev_edge_triggered0_re) begin
        irqarray9_edge_triggered_storage[15:0] <= csrbank22_ev_edge_triggered0_r;
    end
    irqarray9_edge_triggered_re <= csrbank22_ev_edge_triggered0_re;
    if (csrbank22_ev_polarity0_re) begin
        irqarray9_polarity_storage[15:0] <= csrbank22_ev_polarity0_r;
    end
    irqarray9_polarity_re <= csrbank22_ev_polarity0_re;
    irqarray9_status_re <= csrbank22_ev_status_re;
    if (csrbank22_ev_pending_re) begin
        irqarray9_pending_r[15:0] <= csrbank22_ev_pending_r;
    end
    irqarray9_pending_re <= csrbank22_ev_pending_re;
    if (csrbank22_ev_enable0_re) begin
        irqarray9_enable_storage[15:0] <= csrbank22_ev_enable0_r;
    end
    irqarray9_enable_re <= csrbank22_ev_enable0_re;
    interface23_bank_bus_dat_r <= 1'd0;
    if (csrbank23_sel) begin
        case (interface23_bank_bus_adr[9:0])
            1'd0: begin
                interface23_bank_bus_dat_r <= csrbank23_wdata0_w;
            end
            1'd1: begin
                interface23_bank_bus_dat_r <= csrbank23_rdata_w;
            end
            2'd2: begin
                interface23_bank_bus_dat_r <= csrbank23_ev_status_w;
            end
            2'd3: begin
                interface23_bank_bus_dat_r <= csrbank23_ev_pending_w;
            end
            3'd4: begin
                interface23_bank_bus_dat_r <= csrbank23_ev_enable0_w;
            end
            3'd5: begin
                interface23_bank_bus_dat_r <= csrbank23_status_w;
            end
            3'd6: begin
                interface23_bank_bus_dat_r <= csrbank23_control0_w;
            end
            3'd7: begin
                interface23_bank_bus_dat_r <= csrbank23_done0_w;
            end
            4'd8: begin
                interface23_bank_bus_dat_r <= csrbank23_loopback0_w;
            end
        endcase
    end
    if (csrbank23_wdata0_re) begin
        mailbox_wdata_storage[31:0] <= csrbank23_wdata0_r;
    end
    mailbox_wdata_re <= csrbank23_wdata0_re;
    mailbox_rdata_re <= csrbank23_rdata_re;
    mailbox_status_re0 <= csrbank23_ev_status_re;
    if (csrbank23_ev_pending_re) begin
        mailbox_pending_r[3:0] <= csrbank23_ev_pending_r;
    end
    mailbox_pending_re <= csrbank23_ev_pending_re;
    if (csrbank23_ev_enable0_re) begin
        mailbox_enable_storage[3:0] <= csrbank23_ev_enable0_r;
    end
    mailbox_enable_re <= csrbank23_ev_enable0_re;
    mailbox_status_re1 <= csrbank23_status_re;
    if (csrbank23_control0_re) begin
        mailbox_control_storage <= csrbank23_control0_r;
    end
    mailbox_control_re <= csrbank23_control0_re;
    if (csrbank23_done0_re) begin
        mailbox_done_storage <= csrbank23_done0_r;
    end
    mailbox_done_re <= csrbank23_done0_re;
    if (csrbank23_loopback0_re) begin
        mailbox_loopback_storage <= csrbank23_loopback0_r;
    end
    mailbox_loopback_re <= csrbank23_loopback0_re;
    interface24_bank_bus_dat_r <= 1'd0;
    if (csrbank24_sel) begin
        case (interface24_bank_bus_adr[9:0])
            1'd0: begin
                interface24_bank_bus_dat_r <= csrbank24_wdata0_w;
            end
            1'd1: begin
                interface24_bank_bus_dat_r <= csrbank24_rdata_w;
            end
            2'd2: begin
                interface24_bank_bus_dat_r <= csrbank24_status_w;
            end
            2'd3: begin
                interface24_bank_bus_dat_r <= csrbank24_ev_status_w;
            end
            3'd4: begin
                interface24_bank_bus_dat_r <= csrbank24_ev_pending_w;
            end
            3'd5: begin
                interface24_bank_bus_dat_r <= csrbank24_ev_enable0_w;
            end
            3'd6: begin
                interface24_bank_bus_dat_r <= csrbank24_control0_w;
            end
            3'd7: begin
                interface24_bank_bus_dat_r <= csrbank24_done0_w;
            end
        endcase
    end
    if (csrbank24_wdata0_re) begin
        mb_client_wdata_storage[31:0] <= csrbank24_wdata0_r;
    end
    mb_client_wdata_re <= csrbank24_wdata0_re;
    mb_client_rdata_re <= csrbank24_rdata_re;
    mb_client_status_re0 <= csrbank24_status_re;
    mb_client_status_re1 <= csrbank24_ev_status_re;
    if (csrbank24_ev_pending_re) begin
        mb_client_pending_r[3:0] <= csrbank24_ev_pending_r;
    end
    mb_client_pending_re <= csrbank24_ev_pending_re;
    if (csrbank24_ev_enable0_re) begin
        mb_client_enable_storage[3:0] <= csrbank24_ev_enable0_r;
    end
    mb_client_enable_re <= csrbank24_ev_enable0_re;
    if (csrbank24_control0_re) begin
        mb_client_control_storage <= csrbank24_control0_r;
    end
    mb_client_control_re <= csrbank24_control0_re;
    if (csrbank24_done0_re) begin
        mb_client_done_storage <= csrbank24_done0_r;
    end
    mb_client_done_re <= csrbank24_done0_re;
    interface25_bank_bus_dat_r <= 1'd0;
    if (csrbank25_sel) begin
        case (interface25_bank_bus_adr[9:0])
            1'd0: begin
                interface25_bank_bus_dat_r <= csrbank25_pc_w;
            end
        endcase
    end
    re <= csrbank25_pc_re;
    interface26_bank_bus_dat_r <= 1'd0;
    if (csrbank26_sel) begin
        case (interface26_bank_bus_adr[9:0])
            1'd0: begin
                interface26_bank_bus_dat_r <= csrbank26_control0_w;
            end
            1'd1: begin
                interface26_bank_bus_dat_r <= csrbank26_resume_time1_w;
            end
            2'd2: begin
                interface26_bank_bus_dat_r <= csrbank26_resume_time0_w;
            end
            2'd3: begin
                interface26_bank_bus_dat_r <= csrbank26_time1_w;
            end
            3'd4: begin
                interface26_bank_bus_dat_r <= csrbank26_time0_w;
            end
            3'd5: begin
                interface26_bank_bus_dat_r <= csrbank26_status_w;
            end
            3'd6: begin
                interface26_bank_bus_dat_r <= csrbank26_state0_w;
            end
            3'd7: begin
                interface26_bank_bus_dat_r <= csrbank26_interrupt0_w;
            end
            4'd8: begin
                interface26_bank_bus_dat_r <= csrbank26_ev_status_w;
            end
            4'd9: begin
                interface26_bank_bus_dat_r <= csrbank26_ev_pending_w;
            end
            4'd10: begin
                interface26_bank_bus_dat_r <= csrbank26_ev_enable0_w;
            end
        endcase
    end
    if (csrbank26_control0_re) begin
        susres_control_storage[1:0] <= csrbank26_control0_r;
    end
    susres_control_re <= csrbank26_control0_re;
    if (csrbank26_resume_time1_re) begin
        susres_resume_time_storage[63:32] <= csrbank26_resume_time1_r;
    end
    if (csrbank26_resume_time0_re) begin
        susres_resume_time_storage[31:0] <= csrbank26_resume_time0_r;
    end
    susres_resume_time_re <= csrbank26_resume_time0_re;
    susres_time_re <= csrbank26_time0_re;
    susres_status_re0 <= csrbank26_status_re;
    if (csrbank26_state0_re) begin
        susres_state_storage[1:0] <= csrbank26_state0_r;
    end
    susres_state_re <= csrbank26_state0_re;
    if (csrbank26_interrupt0_re) begin
        susres_interrupt_storage <= csrbank26_interrupt0_r;
    end
    susres_interrupt_re <= csrbank26_interrupt0_re;
    susres_status_re1 <= csrbank26_ev_status_re;
    if (csrbank26_ev_pending_re) begin
        susres_pending_r <= csrbank26_ev_pending_r;
    end
    susres_pending_re <= csrbank26_ev_pending_re;
    if (csrbank26_ev_enable0_re) begin
        susres_enable_storage <= csrbank26_ev_enable0_r;
    end
    susres_enable_re <= csrbank26_ev_enable0_re;
    interface27_bank_bus_dat_r <= 1'd0;
    if (csrbank27_sel) begin
        case (interface27_bank_bus_adr[9:0])
            1'd0: begin
                interface27_bank_bus_dat_r <= csrbank27_control0_w;
            end
            1'd1: begin
                interface27_bank_bus_dat_r <= csrbank27_time1_w;
            end
            2'd2: begin
                interface27_bank_bus_dat_r <= csrbank27_time0_w;
            end
            2'd3: begin
                interface27_bank_bus_dat_r <= csrbank27_msleep_target1_w;
            end
            3'd4: begin
                interface27_bank_bus_dat_r <= csrbank27_msleep_target0_w;
            end
            3'd5: begin
                interface27_bank_bus_dat_r <= csrbank27_ev_status_w;
            end
            3'd6: begin
                interface27_bank_bus_dat_r <= csrbank27_ev_pending_w;
            end
            3'd7: begin
                interface27_bank_bus_dat_r <= csrbank27_ev_enable0_w;
            end
            4'd8: begin
                interface27_bank_bus_dat_r <= csrbank27_clocks_per_tick0_w;
            end
        endcase
    end
    if (csrbank27_control0_re) begin
        ticktimer_control_storage <= csrbank27_control0_r;
    end
    ticktimer_control_re <= csrbank27_control0_re;
    ticktimer_time_re <= csrbank27_time0_re;
    if (csrbank27_msleep_target1_re) begin
        ticktimer_msleep_target_storage[63:32] <= csrbank27_msleep_target1_r;
    end
    if (csrbank27_msleep_target0_re) begin
        ticktimer_msleep_target_storage[31:0] <= csrbank27_msleep_target0_r;
    end
    ticktimer_msleep_target_re <= csrbank27_msleep_target0_re;
    ticktimer_status_re <= csrbank27_ev_status_re;
    if (csrbank27_ev_pending_re) begin
        ticktimer_pending_r <= csrbank27_ev_pending_r;
    end
    ticktimer_pending_re <= csrbank27_ev_pending_re;
    if (csrbank27_ev_enable0_re) begin
        ticktimer_enable_storage <= csrbank27_ev_enable0_r;
    end
    ticktimer_enable_re <= csrbank27_ev_enable0_re;
    if (csrbank27_clocks_per_tick0_re) begin
        ticktimer_clocks_per_tick_storage[31:0] <= csrbank27_clocks_per_tick0_r;
    end
    ticktimer_clocks_per_tick_re <= csrbank27_clocks_per_tick0_re;
    interface28_bank_bus_dat_r <= 1'd0;
    if (csrbank28_sel) begin
        case (interface28_bank_bus_adr[9:0])
            1'd0: begin
                interface28_bank_bus_dat_r <= csrbank28_load0_w;
            end
            1'd1: begin
                interface28_bank_bus_dat_r <= csrbank28_reload0_w;
            end
            2'd2: begin
                interface28_bank_bus_dat_r <= csrbank28_en0_w;
            end
            2'd3: begin
                interface28_bank_bus_dat_r <= csrbank28_update_value0_w;
            end
            3'd4: begin
                interface28_bank_bus_dat_r <= csrbank28_value_w;
            end
            3'd5: begin
                interface28_bank_bus_dat_r <= csrbank28_ev_status_w;
            end
            3'd6: begin
                interface28_bank_bus_dat_r <= csrbank28_ev_pending_w;
            end
            3'd7: begin
                interface28_bank_bus_dat_r <= csrbank28_ev_enable0_w;
            end
        endcase
    end
    if (csrbank28_load0_re) begin
        cramsoc_load_storage[31:0] <= csrbank28_load0_r;
    end
    cramsoc_load_re <= csrbank28_load0_re;
    if (csrbank28_reload0_re) begin
        cramsoc_reload_storage[31:0] <= csrbank28_reload0_r;
    end
    cramsoc_reload_re <= csrbank28_reload0_re;
    if (csrbank28_en0_re) begin
        cramsoc_en_storage <= csrbank28_en0_r;
    end
    cramsoc_en_re <= csrbank28_en0_re;
    if (csrbank28_update_value0_re) begin
        cramsoc_update_value_storage <= csrbank28_update_value0_r;
    end
    cramsoc_update_value_re <= csrbank28_update_value0_re;
    cramsoc_value_re <= csrbank28_value_re;
    cramsoc_status_re <= csrbank28_ev_status_re;
    if (csrbank28_ev_pending_re) begin
        cramsoc_pending_r <= csrbank28_ev_pending_r;
    end
    cramsoc_pending_re <= csrbank28_ev_pending_re;
    if (csrbank28_ev_enable0_re) begin
        cramsoc_enable_storage <= csrbank28_ev_enable0_r;
    end
    cramsoc_enable_re <= csrbank28_ev_enable0_re;
    if (sys_rst) begin
        cramsoc_load_storage <= 32'd0;
        cramsoc_load_re <= 1'd0;
        cramsoc_reload_storage <= 32'd0;
        cramsoc_reload_re <= 1'd0;
        cramsoc_en_storage <= 1'd0;
        cramsoc_en_re <= 1'd0;
        cramsoc_update_value_storage <= 1'd0;
        cramsoc_update_value_re <= 1'd0;
        cramsoc_value_status <= 32'd0;
        cramsoc_value_re <= 1'd0;
        cramsoc_zero_pending <= 1'd0;
        cramsoc_zero_trigger_d <= 1'd0;
        cramsoc_status_re <= 1'd0;
        cramsoc_pending_re <= 1'd0;
        cramsoc_pending_r <= 1'd0;
        cramsoc_enable_storage <= 1'd0;
        cramsoc_enable_re <= 1'd0;
        cramsoc_value <= 32'd0;
        reset_debug_logic <= 1'd0;
        debug_reset <= 1'd0;
        re <= 1'd0;
        coreuser_vex <= 8'd0;
        vex_mm <= 1'd0;
        coreuser_control_storage <= 2'd0;
        coreuser_control_re <= 1'd0;
        coreuser_coreuser <= 8'd0;
        coreuser_mm <= 1'd0;
        coreuser_status_re <= 1'd0;
        coreuser_map_lo_storage <= 32'd0;
        coreuser_map_lo_re <= 1'd0;
        coreuser_map_hi_storage <= 32'd0;
        coreuser_map_hi_re <= 1'd0;
        coreuser_uservalue_storage <= 18'd0;
        coreuser_uservalue_re <= 1'd0;
        coreuser_protect_storage <= 1'd0;
        coreuser_protect_re <= 1'd0;
        coreuser_enable1 <= 1'd0;
        coreuser_invert_priv1 <= 1'd0;
        coreuser_lut01 <= 8'd0;
        coreuser_lut11 <= 8'd0;
        coreuser_lut21 <= 8'd0;
        coreuser_lut31 <= 8'd0;
        coreuser_lut41 <= 8'd0;
        coreuser_lut51 <= 8'd0;
        coreuser_lut61 <= 8'd0;
        coreuser_lut71 <= 8'd0;
        coreuser_user01 <= 2'd0;
        coreuser_user11 <= 2'd0;
        coreuser_user21 <= 2'd0;
        coreuser_user31 <= 2'd0;
        coreuser_user41 <= 2'd0;
        coreuser_user51 <= 2'd0;
        coreuser_user61 <= 2'd0;
        coreuser_user71 <= 2'd0;
        coreuser_user_default <= 2'd0;
        ibus_r_active <= 1'd0;
        dbus_r_active <= 1'd0;
        dbus_w_active <= 1'd0;
        pbus_r_active <= 1'd0;
        pbus_w_active <= 1'd0;
        active_timeout <= 7'd0;
        irqarray0_soft_storage <= 16'd0;
        irqarray0_soft_re <= 1'd0;
        irqarray0_edge_triggered_storage <= 16'd0;
        irqarray0_edge_triggered_re <= 1'd0;
        irqarray0_polarity_storage <= 16'd0;
        irqarray0_polarity_re <= 1'd0;
        irqarray0_status_re <= 1'd0;
        irqarray0_pending_re <= 1'd0;
        irqarray0_pending_r <= 16'd0;
        irqarray0_enable_storage <= 16'd0;
        irqarray0_enable_re <= 1'd0;
        irqarray1_soft_storage <= 16'd0;
        irqarray1_soft_re <= 1'd0;
        irqarray1_edge_triggered_storage <= 16'd0;
        irqarray1_edge_triggered_re <= 1'd0;
        irqarray1_polarity_storage <= 16'd0;
        irqarray1_polarity_re <= 1'd0;
        irqarray1_status_re <= 1'd0;
        irqarray1_pending_re <= 1'd0;
        irqarray1_pending_r <= 16'd0;
        irqarray1_enable_storage <= 16'd0;
        irqarray1_enable_re <= 1'd0;
        irqarray2_soft_storage <= 16'd0;
        irqarray2_soft_re <= 1'd0;
        irqarray2_edge_triggered_storage <= 16'd0;
        irqarray2_edge_triggered_re <= 1'd0;
        irqarray2_polarity_storage <= 16'd0;
        irqarray2_polarity_re <= 1'd0;
        irqarray2_status_re <= 1'd0;
        irqarray2_pending_re <= 1'd0;
        irqarray2_pending_r <= 16'd0;
        irqarray2_enable_storage <= 16'd0;
        irqarray2_enable_re <= 1'd0;
        irqarray3_soft_storage <= 16'd0;
        irqarray3_soft_re <= 1'd0;
        irqarray3_edge_triggered_storage <= 16'd0;
        irqarray3_edge_triggered_re <= 1'd0;
        irqarray3_polarity_storage <= 16'd0;
        irqarray3_polarity_re <= 1'd0;
        irqarray3_status_re <= 1'd0;
        irqarray3_pending_re <= 1'd0;
        irqarray3_pending_r <= 16'd0;
        irqarray3_enable_storage <= 16'd0;
        irqarray3_enable_re <= 1'd0;
        irqarray4_soft_storage <= 16'd0;
        irqarray4_soft_re <= 1'd0;
        irqarray4_edge_triggered_storage <= 16'd0;
        irqarray4_edge_triggered_re <= 1'd0;
        irqarray4_polarity_storage <= 16'd0;
        irqarray4_polarity_re <= 1'd0;
        irqarray4_status_re <= 1'd0;
        irqarray4_pending_re <= 1'd0;
        irqarray4_pending_r <= 16'd0;
        irqarray4_enable_storage <= 16'd0;
        irqarray4_enable_re <= 1'd0;
        irqarray5_soft_storage <= 16'd0;
        irqarray5_soft_re <= 1'd0;
        irqarray5_edge_triggered_storage <= 16'd0;
        irqarray5_edge_triggered_re <= 1'd0;
        irqarray5_polarity_storage <= 16'd0;
        irqarray5_polarity_re <= 1'd0;
        irqarray5_status_re <= 1'd0;
        irqarray5_pending_re <= 1'd0;
        irqarray5_pending_r <= 16'd0;
        irqarray5_enable_storage <= 16'd0;
        irqarray5_enable_re <= 1'd0;
        irqarray6_soft_storage <= 16'd0;
        irqarray6_soft_re <= 1'd0;
        irqarray6_edge_triggered_storage <= 16'd0;
        irqarray6_edge_triggered_re <= 1'd0;
        irqarray6_polarity_storage <= 16'd0;
        irqarray6_polarity_re <= 1'd0;
        irqarray6_status_re <= 1'd0;
        irqarray6_pending_re <= 1'd0;
        irqarray6_pending_r <= 16'd0;
        irqarray6_enable_storage <= 16'd0;
        irqarray6_enable_re <= 1'd0;
        irqarray7_soft_storage <= 16'd0;
        irqarray7_soft_re <= 1'd0;
        irqarray7_edge_triggered_storage <= 16'd0;
        irqarray7_edge_triggered_re <= 1'd0;
        irqarray7_polarity_storage <= 16'd0;
        irqarray7_polarity_re <= 1'd0;
        irqarray7_status_re <= 1'd0;
        irqarray7_pending_re <= 1'd0;
        irqarray7_pending_r <= 16'd0;
        irqarray7_enable_storage <= 16'd0;
        irqarray7_enable_re <= 1'd0;
        irqarray8_soft_storage <= 16'd0;
        irqarray8_soft_re <= 1'd0;
        irqarray8_edge_triggered_storage <= 16'd0;
        irqarray8_edge_triggered_re <= 1'd0;
        irqarray8_polarity_storage <= 16'd0;
        irqarray8_polarity_re <= 1'd0;
        irqarray8_status_re <= 1'd0;
        irqarray8_pending_re <= 1'd0;
        irqarray8_pending_r <= 16'd0;
        irqarray8_enable_storage <= 16'd0;
        irqarray8_enable_re <= 1'd0;
        irqarray9_soft_storage <= 16'd0;
        irqarray9_soft_re <= 1'd0;
        irqarray9_edge_triggered_storage <= 16'd0;
        irqarray9_edge_triggered_re <= 1'd0;
        irqarray9_polarity_storage <= 16'd0;
        irqarray9_polarity_re <= 1'd0;
        irqarray9_status_re <= 1'd0;
        irqarray9_pending_re <= 1'd0;
        irqarray9_pending_r <= 16'd0;
        irqarray9_enable_storage <= 16'd0;
        irqarray9_enable_re <= 1'd0;
        irqarray10_soft_storage <= 16'd0;
        irqarray10_soft_re <= 1'd0;
        irqarray10_edge_triggered_storage <= 16'd0;
        irqarray10_edge_triggered_re <= 1'd0;
        irqarray10_polarity_storage <= 16'd0;
        irqarray10_polarity_re <= 1'd0;
        irqarray10_status_re <= 1'd0;
        irqarray10_pending_re <= 1'd0;
        irqarray10_pending_r <= 16'd0;
        irqarray10_enable_storage <= 16'd0;
        irqarray10_enable_re <= 1'd0;
        irqarray11_soft_storage <= 16'd0;
        irqarray11_soft_re <= 1'd0;
        irqarray11_edge_triggered_storage <= 16'd0;
        irqarray11_edge_triggered_re <= 1'd0;
        irqarray11_polarity_storage <= 16'd0;
        irqarray11_polarity_re <= 1'd0;
        irqarray11_status_re <= 1'd0;
        irqarray11_pending_re <= 1'd0;
        irqarray11_pending_r <= 16'd0;
        irqarray11_enable_storage <= 16'd0;
        irqarray11_enable_re <= 1'd0;
        irqarray12_soft_storage <= 16'd0;
        irqarray12_soft_re <= 1'd0;
        irqarray12_edge_triggered_storage <= 16'd0;
        irqarray12_edge_triggered_re <= 1'd0;
        irqarray12_polarity_storage <= 16'd0;
        irqarray12_polarity_re <= 1'd0;
        irqarray12_status_re <= 1'd0;
        irqarray12_pending_re <= 1'd0;
        irqarray12_pending_r <= 16'd0;
        irqarray12_enable_storage <= 16'd0;
        irqarray12_enable_re <= 1'd0;
        irqarray13_soft_storage <= 16'd0;
        irqarray13_soft_re <= 1'd0;
        irqarray13_edge_triggered_storage <= 16'd0;
        irqarray13_edge_triggered_re <= 1'd0;
        irqarray13_polarity_storage <= 16'd0;
        irqarray13_polarity_re <= 1'd0;
        irqarray13_status_re <= 1'd0;
        irqarray13_pending_re <= 1'd0;
        irqarray13_pending_r <= 16'd0;
        irqarray13_enable_storage <= 16'd0;
        irqarray13_enable_re <= 1'd0;
        irqarray14_soft_storage <= 16'd0;
        irqarray14_soft_re <= 1'd0;
        irqarray14_edge_triggered_storage <= 16'd0;
        irqarray14_edge_triggered_re <= 1'd0;
        irqarray14_polarity_storage <= 16'd0;
        irqarray14_polarity_re <= 1'd0;
        irqarray14_status_re <= 1'd0;
        irqarray14_pending_re <= 1'd0;
        irqarray14_pending_r <= 16'd0;
        irqarray14_enable_storage <= 16'd0;
        irqarray14_enable_re <= 1'd0;
        irqarray15_soft_storage <= 16'd0;
        irqarray15_soft_re <= 1'd0;
        irqarray15_edge_triggered_storage <= 16'd0;
        irqarray15_edge_triggered_re <= 1'd0;
        irqarray15_polarity_storage <= 16'd0;
        irqarray15_polarity_re <= 1'd0;
        irqarray15_status_re <= 1'd0;
        irqarray15_pending_re <= 1'd0;
        irqarray15_pending_r <= 16'd0;
        irqarray15_enable_storage <= 16'd0;
        irqarray15_enable_re <= 1'd0;
        irqarray16_soft_storage <= 16'd0;
        irqarray16_soft_re <= 1'd0;
        irqarray16_edge_triggered_storage <= 16'd0;
        irqarray16_edge_triggered_re <= 1'd0;
        irqarray16_polarity_storage <= 16'd0;
        irqarray16_polarity_re <= 1'd0;
        irqarray16_status_re <= 1'd0;
        irqarray16_pending_re <= 1'd0;
        irqarray16_pending_r <= 16'd0;
        irqarray16_enable_storage <= 16'd0;
        irqarray16_enable_re <= 1'd0;
        irqarray17_soft_storage <= 16'd0;
        irqarray17_soft_re <= 1'd0;
        irqarray17_edge_triggered_storage <= 16'd0;
        irqarray17_edge_triggered_re <= 1'd0;
        irqarray17_polarity_storage <= 16'd0;
        irqarray17_polarity_re <= 1'd0;
        irqarray17_status_re <= 1'd0;
        irqarray17_pending_re <= 1'd0;
        irqarray17_pending_r <= 16'd0;
        irqarray17_enable_storage <= 16'd0;
        irqarray17_enable_re <= 1'd0;
        irqarray18_soft_storage <= 16'd0;
        irqarray18_soft_re <= 1'd0;
        irqarray18_edge_triggered_storage <= 16'd0;
        irqarray18_edge_triggered_re <= 1'd0;
        irqarray18_polarity_storage <= 16'd0;
        irqarray18_polarity_re <= 1'd0;
        irqarray18_status_re <= 1'd0;
        irqarray18_pending_re <= 1'd0;
        irqarray18_pending_r <= 16'd0;
        irqarray18_enable_storage <= 16'd0;
        irqarray18_enable_re <= 1'd0;
        irqarray19_soft_storage <= 16'd0;
        irqarray19_soft_re <= 1'd0;
        irqarray19_edge_triggered_storage <= 16'd0;
        irqarray19_edge_triggered_re <= 1'd0;
        irqarray19_polarity_storage <= 16'd0;
        irqarray19_polarity_re <= 1'd0;
        irqarray19_status_re <= 1'd0;
        irqarray19_pending_re <= 1'd0;
        irqarray19_pending_r <= 16'd0;
        irqarray19_enable_storage <= 16'd0;
        irqarray19_enable_re <= 1'd0;
        ticktimer_control_storage <= 1'd0;
        ticktimer_control_re <= 1'd0;
        ticktimer_time_re <= 1'd0;
        ticktimer_msleep_target_storage <= 64'd0;
        ticktimer_msleep_target_re <= 1'd0;
        ticktimer_status_re <= 1'd0;
        ticktimer_pending_re <= 1'd0;
        ticktimer_pending_r <= 1'd0;
        ticktimer_enable_storage <= 1'd0;
        ticktimer_enable_re <= 1'd0;
        ticktimer_clocks_per_tick_storage <= 32'd800000;
        ticktimer_clocks_per_tick_re <= 1'd0;
        d11ctime_control_storage <= 32'd400000;
        d11ctime_control_re <= 1'd0;
        d11ctime_heartbeat_re <= 1'd0;
        susres_control_storage <= 2'd0;
        susres_control_re <= 1'd0;
        susres_resume_time_storage <= 64'd0;
        susres_resume_time_re <= 1'd0;
        susres_time_re <= 1'd0;
        susres_status_re0 <= 1'd0;
        susres_state_storage <= 2'd0;
        susres_state_re <= 1'd0;
        susres_interrupt_storage <= 1'd0;
        susres_interrupt_re <= 1'd0;
        susres_status_re1 <= 1'd0;
        susres_pending_re <= 1'd0;
        susres_pending_r <= 1'd0;
        susres_enable_storage <= 1'd0;
        susres_enable_re <= 1'd0;
        mailbox_w_abort <= 1'd0;
        mailbox_wdata_storage <= 32'd0;
        mailbox_wdata_re <= 1'd0;
        mailbox_rdata_re <= 1'd0;
        mailbox_available_pending <= 1'd0;
        mailbox_abort_init_pending <= 1'd0;
        mailbox_abort_init_trigger_d <= 1'd0;
        mailbox_abort_done_pending <= 1'd0;
        mailbox_abort_done_trigger_d <= 1'd0;
        mailbox_error_pending <= 1'd0;
        mailbox_error_trigger_d <= 1'd0;
        mailbox_status_re0 <= 1'd0;
        mailbox_pending_re <= 1'd0;
        mailbox_pending_r <= 4'd0;
        mailbox_enable_storage <= 4'd0;
        mailbox_enable_re <= 1'd0;
        mailbox_status_re1 <= 1'd0;
        mailbox_control_storage <= 1'd0;
        mailbox_control_re <= 1'd0;
        mailbox_done_storage <= 1'd0;
        mailbox_done_re <= 1'd0;
        mailbox_loopback_storage <= 1'd0;
        mailbox_loopback_re <= 1'd0;
        mailbox_abort_in_progress1 <= 1'd0;
        mailbox_abort_ack1 <= 1'd0;
        mailbox_w_over_bit <= 1'd0;
        mailbox_syncfifobufferedmacro0_syncfifobufferedmacro0_readable <= 1'd0;
        mailbox_syncfifobufferedmacro0_fifo_level <= 11'd0;
        mailbox_syncfifobufferedmacro0_fifo_produce <= 10'd0;
        mailbox_syncfifobufferedmacro0_fifo_consume <= 10'd0;
        mailbox_r_over_bit <= 1'd0;
        mailbox_syncfifobufferedmacro1_syncfifobufferedmacro1_readable <= 1'd0;
        mailbox_syncfifobufferedmacro1_fifo_level <= 11'd0;
        mailbox_syncfifobufferedmacro1_fifo_produce <= 10'd0;
        mailbox_syncfifobufferedmacro1_fifo_consume <= 10'd0;
        mb_client_w_abort <= 1'd0;
        mb_client_wdata_storage <= 32'd0;
        mb_client_wdata_re <= 1'd0;
        mb_client_rdata_re <= 1'd0;
        mb_client_tx_err <= 1'd0;
        mb_client_rx_err <= 1'd0;
        mb_client_status_re0 <= 1'd0;
        mb_client_available_pending <= 1'd0;
        mb_client_abort_init_pending <= 1'd0;
        mb_client_abort_init_trigger_d <= 1'd0;
        mb_client_abort_done_pending <= 1'd0;
        mb_client_abort_done_trigger_d <= 1'd0;
        mb_client_error_pending <= 1'd0;
        mb_client_error_trigger_d <= 1'd0;
        mb_client_status_re1 <= 1'd0;
        mb_client_pending_re <= 1'd0;
        mb_client_pending_r <= 4'd0;
        mb_client_enable_storage <= 4'd0;
        mb_client_enable_re <= 1'd0;
        mb_client_control_storage <= 1'd0;
        mb_client_control_re <= 1'd0;
        mb_client_done_storage <= 1'd0;
        mb_client_done_re <= 1'd0;
        mb_client_abort_in_progress1 <= 1'd0;
        mb_client_abort_ack1 <= 1'd0;
        mb_client_w_pending <= 1'd0;
        csr_wtest_storage <= 32'd0;
        csr_wtest_re <= 1'd0;
        csr_rtest_re <= 1'd0;
        cramsoc_last_was_read <= 1'd0;
        socbushandler_slave_sel_reg0 <= 1'd0;
        socbushandler_slave_sel_reg1 <= 1'd0;
        socbushandler_axiliterequestcounter0_counter <= 8'd0;
        socbushandler_axiliterequestcounter1_counter <= 8'd0;
        socbushandler_wr_lock_counter <= 8'd0;
        socbushandler_rd_lock_counter <= 8'd0;
        cramsoc_mailbox_state <= 2'd0;
        cramsoc_mailboxclient_state <= 2'd0;
        cramsoc_axilite2csr_state <= 2'd0;
    end
end


//------------------------------------------------------------------------------
// Specialized Logic
//------------------------------------------------------------------------------

axi_axil_adapter #(
	.ADDR_WIDTH(6'd32),
	.AXIL_DATA_WIDTH(6'd32),
	.AXI_DATA_WIDTH(6'd32),
	.AXI_ID_WIDTH(1'd1),
	.CONVERT_BURST(1'd1),
	.CONVERT_NARROW_BURST(1'd0)
) axi_axil_adapter (
	.clk(sys_clk),
	.m_axil_arready(cramsoc_peripherals_ar_ready),
	.m_axil_awready(cramsoc_peripherals_aw_ready),
	.m_axil_bresp(cramsoc_peripherals_b_payload_resp),
	.m_axil_bvalid(cramsoc_peripherals_b_valid),
	.m_axil_rdata(cramsoc_peripherals_r_payload_data),
	.m_axil_rresp(cramsoc_peripherals_r_payload_resp),
	.m_axil_rvalid(cramsoc_peripherals_r_valid),
	.m_axil_wready(cramsoc_peripherals_w_ready),
	.rst(sys_rst),
	.s_axi_araddr(cramsoc_dbus_peri_ar_payload_addr),
	.s_axi_arburst(cramsoc_dbus_peri_ar_payload_burst),
	.s_axi_arcache(cramsoc_dbus_peri_ar_payload_cache),
	.s_axi_arid(cramsoc_dbus_peri_ar_param_id),
	.s_axi_arlen(cramsoc_dbus_peri_ar_payload_len),
	.s_axi_arlock(cramsoc_dbus_peri_ar_payload_lock),
	.s_axi_arprot(cramsoc_dbus_peri_ar_payload_prot),
	.s_axi_arsize(cramsoc_dbus_peri_ar_payload_size),
	.s_axi_arvalid(cramsoc_dbus_peri_ar_valid),
	.s_axi_awaddr(cramsoc_dbus_peri_aw_payload_addr),
	.s_axi_awburst(cramsoc_dbus_peri_aw_payload_burst),
	.s_axi_awcache(cramsoc_dbus_peri_aw_payload_cache),
	.s_axi_awid(cramsoc_dbus_peri_aw_param_id),
	.s_axi_awlen(cramsoc_dbus_peri_aw_payload_len),
	.s_axi_awlock(cramsoc_dbus_peri_aw_payload_lock),
	.s_axi_awprot(cramsoc_dbus_peri_aw_payload_prot),
	.s_axi_awsize(cramsoc_dbus_peri_aw_payload_size),
	.s_axi_awvalid(cramsoc_dbus_peri_aw_valid),
	.s_axi_bready(cramsoc_dbus_peri_b_ready),
	.s_axi_rready(cramsoc_dbus_peri_r_ready),
	.s_axi_wdata(cramsoc_dbus_peri_w_payload_data),
	.s_axi_wlast(cramsoc_dbus_peri_w_last),
	.s_axi_wstrb(cramsoc_dbus_peri_w_payload_strb),
	.s_axi_wvalid(cramsoc_dbus_peri_w_valid),
	.m_axil_araddr(cramsoc_peripherals_ar_payload_addr),
	.m_axil_arprot(cramsoc_peripherals_ar_payload_prot),
	.m_axil_arvalid(cramsoc_peripherals_ar_valid),
	.m_axil_awaddr(cramsoc_peripherals_aw_payload_addr),
	.m_axil_awprot(cramsoc_peripherals_aw_payload_prot),
	.m_axil_awvalid(cramsoc_peripherals_aw_valid),
	.m_axil_bready(cramsoc_peripherals_b_ready),
	.m_axil_rready(cramsoc_peripherals_r_ready),
	.m_axil_wdata(cramsoc_peripherals_w_payload_data),
	.m_axil_wstrb(cramsoc_peripherals_w_payload_strb),
	.m_axil_wvalid(cramsoc_peripherals_w_valid),
	.s_axi_arready(cramsoc_dbus_peri_ar_ready),
	.s_axi_awready(cramsoc_dbus_peri_aw_ready),
	.s_axi_bid(cramsoc_dbus_peri_b_param_id),
	.s_axi_bresp(cramsoc_dbus_peri_b_payload_resp),
	.s_axi_bvalid(cramsoc_dbus_peri_b_valid),
	.s_axi_rdata(cramsoc_dbus_peri_r_payload_data),
	.s_axi_rid(cramsoc_dbus_peri_r_param_id),
	.s_axi_rlast(cramsoc_dbus_peri_r_last),
	.s_axi_rresp(cramsoc_dbus_peri_r_payload_resp),
	.s_axi_rvalid(cramsoc_dbus_peri_r_valid),
	.s_axi_wready(cramsoc_dbus_peri_w_ready)
);

axi_axil_adapter #(
	.ADDR_WIDTH(6'd32),
	.AXIL_DATA_WIDTH(6'd32),
	.AXI_DATA_WIDTH(6'd32),
	.AXI_ID_WIDTH(1'd1),
	.CONVERT_BURST(1'd1),
	.CONVERT_NARROW_BURST(1'd0)
) axi_axil_adapter_1 (
	.clk(sys_clk),
	.m_axil_arready(cramsoc_corecsr_ar_ready),
	.m_axil_awready(cramsoc_corecsr_aw_ready),
	.m_axil_bresp(cramsoc_corecsr_b_payload_resp),
	.m_axil_bvalid(cramsoc_corecsr_b_valid),
	.m_axil_rdata(cramsoc_corecsr_r_payload_data),
	.m_axil_rresp(cramsoc_corecsr_r_payload_resp),
	.m_axil_rvalid(cramsoc_corecsr_r_valid),
	.m_axil_wready(cramsoc_corecsr_w_ready),
	.rst(sys_rst),
	.s_axi_araddr(cramsoc_axi_csr_ar_payload_addr),
	.s_axi_arburst(cramsoc_axi_csr_ar_payload_burst),
	.s_axi_arcache(cramsoc_axi_csr_ar_payload_cache),
	.s_axi_arid(cramsoc_axi_csr_ar_param_id),
	.s_axi_arlen(cramsoc_axi_csr_ar_payload_len),
	.s_axi_arlock(cramsoc_axi_csr_ar_payload_lock),
	.s_axi_arprot(cramsoc_axi_csr_ar_payload_prot),
	.s_axi_arsize(cramsoc_axi_csr_ar_payload_size),
	.s_axi_arvalid(cramsoc_axi_csr_ar_valid),
	.s_axi_awaddr(cramsoc_axi_csr_aw_payload_addr),
	.s_axi_awburst(cramsoc_axi_csr_aw_payload_burst),
	.s_axi_awcache(cramsoc_axi_csr_aw_payload_cache),
	.s_axi_awid(cramsoc_axi_csr_aw_param_id),
	.s_axi_awlen(cramsoc_axi_csr_aw_payload_len),
	.s_axi_awlock(cramsoc_axi_csr_aw_payload_lock),
	.s_axi_awprot(cramsoc_axi_csr_aw_payload_prot),
	.s_axi_awsize(cramsoc_axi_csr_aw_payload_size),
	.s_axi_awvalid(cramsoc_axi_csr_aw_valid),
	.s_axi_bready(cramsoc_axi_csr_b_ready),
	.s_axi_rready(cramsoc_axi_csr_r_ready),
	.s_axi_wdata(cramsoc_axi_csr_w_payload_data),
	.s_axi_wlast(cramsoc_axi_csr_w_last),
	.s_axi_wstrb(cramsoc_axi_csr_w_payload_strb),
	.s_axi_wvalid(cramsoc_axi_csr_w_valid),
	.m_axil_araddr(cramsoc_corecsr_ar_payload_addr),
	.m_axil_arprot(cramsoc_corecsr_ar_payload_prot),
	.m_axil_arvalid(cramsoc_corecsr_ar_valid),
	.m_axil_awaddr(cramsoc_corecsr_aw_payload_addr),
	.m_axil_awprot(cramsoc_corecsr_aw_payload_prot),
	.m_axil_awvalid(cramsoc_corecsr_aw_valid),
	.m_axil_bready(cramsoc_corecsr_b_ready),
	.m_axil_rready(cramsoc_corecsr_r_ready),
	.m_axil_wdata(cramsoc_corecsr_w_payload_data),
	.m_axil_wstrb(cramsoc_corecsr_w_payload_strb),
	.m_axil_wvalid(cramsoc_corecsr_w_valid),
	.s_axi_arready(cramsoc_axi_csr_ar_ready),
	.s_axi_awready(cramsoc_axi_csr_aw_ready),
	.s_axi_bid(cramsoc_axi_csr_b_param_id),
	.s_axi_bresp(cramsoc_axi_csr_b_payload_resp),
	.s_axi_bvalid(cramsoc_axi_csr_b_valid),
	.s_axi_rdata(cramsoc_axi_csr_r_payload_data),
	.s_axi_rid(cramsoc_axi_csr_r_param_id),
	.s_axi_rlast(cramsoc_axi_csr_r_last),
	.s_axi_rresp(cramsoc_axi_csr_r_payload_resp),
	.s_axi_rvalid(cramsoc_axi_csr_r_valid),
	.s_axi_wready(cramsoc_axi_csr_w_ready)
);

fdre_cosim fdre_cosim(
	.C(sys_clk),
	.CE(coreuser_protect_storage),
	.D(1'd1),
	.R(sys_rst),
	.Q(coreuser_protect)
);

Ram_1w_1rs #(
	.clockCrossing(1'd0),
	.ramname("RAM_DP_1024_32"),
	.rdAddressWidth(4'd10),
	.rdDataWidth(6'd32),
	.wordCount(11'd1024),
	.wordWidth(6'd32),
	.wrAddressWidth(4'd10),
	.wrDataWidth(6'd32),
	.wrMaskEnable(1'd0)
) Ram_1w_1rs (
		.rbs	(rbif_rdram1kx32[0]),
	.CMATPG(mailbox_syncfifobufferedmacro0_fifo_cmatpg),
	.CMBIST(mailbox_syncfifobufferedmacro0_fifo_cmbist),
	.rd_addr(mailbox_syncfifobufferedmacro0_fifo_rdport_adr),
	.rd_clk(sys_clk),
	.rd_en(mailbox_syncfifobufferedmacro0_fifo_rdport_re),
	.sramtrm(mailbox_syncfifobufferedmacro0_fifo_vexsramtrm),
	.wr_addr(mailbox_syncfifobufferedmacro0_fifo_wrport_adr),
	.wr_clk(sys_clk),
	.wr_data(mailbox_syncfifobufferedmacro0_fifo_wrport_dat_w),
	.wr_en(mailbox_syncfifobufferedmacro0_fifo_wrport_we),
	.wr_mask(1'd0),
	.rd_data(mailbox_syncfifobufferedmacro0_fifo_rdport_dat_r)
);

Ram_1w_1rs #(
	.clockCrossing(1'd0),
	.ramname("RAM_DP_1024_32"),
	.rdAddressWidth(4'd10),
	.rdDataWidth(6'd32),
	.wordCount(11'd1024),
	.wordWidth(6'd32),
	.wrAddressWidth(4'd10),
	.wrDataWidth(6'd32),
	.wrMaskEnable(1'd0)
) Ram_1w_1rs_1 (
		.rbs	(rbif_rdram1kx32[1]),
	.CMATPG(mailbox_syncfifobufferedmacro1_fifo_cmatpg),
	.CMBIST(mailbox_syncfifobufferedmacro1_fifo_cmbist),
	.rd_addr(mailbox_syncfifobufferedmacro1_fifo_rdport_adr),
	.rd_clk(sys_clk),
	.rd_en(mailbox_syncfifobufferedmacro1_fifo_rdport_re),
	.sramtrm(mailbox_syncfifobufferedmacro1_fifo_vexsramtrm),
	.wr_addr(mailbox_syncfifobufferedmacro1_fifo_wrport_adr),
	.wr_clk(sys_clk),
	.wr_data(mailbox_syncfifobufferedmacro1_fifo_wrport_dat_w),
	.wr_en(mailbox_syncfifobufferedmacro1_fifo_wrport_we),
	.wr_mask(1'd0),
	.rd_data(mailbox_syncfifobufferedmacro1_fifo_rdport_dat_r)
);

axi_crossbar #(
	.ADDR_WIDTH(6'd32),
	.ARUSER_ENABLE(1'd0),
	.ARUSER_WIDTH(1'd1),
	.AWUSER_ENABLE(1'd0),
	.AWUSER_WIDTH(1'd1),
	.BUSER_ENABLE(1'd0),
	.BUSER_WIDTH(1'd1),
	.DATA_WIDTH(6'd32),
	.M_ADDR_WIDTH(96'd534955578257836081181),
	.M_AR_REG_TYPE(6'd21),
	.M_AW_REG_TYPE(6'd21),
	.M_BASE_ADDR(96'd29710560958990027663148580864),
	.M_B_REG_TYPE(6'd21),
	.M_COUNT(2'd3),
	.M_ID_WIDTH(1'd1),
	.M_R_REG_TYPE(6'd42),
	.M_W_REG_TYPE(6'd42),
	.RUSER_ENABLE(1'd0),
	.RUSER_WIDTH(1'd1),
	.S_AR_REG_TYPE(2'd0),
	.S_AW_REG_TYPE(2'd0),
	.S_B_REG_TYPE(2'd0),
	.S_COUNT(1'd1),
	.S_ID_WIDTH(1'd1),
	.S_R_REG_TYPE(2'd0),
	.S_W_REG_TYPE(2'd0),
	.WUSER_ENABLE(1'd0),
	.WUSER_WIDTH(1'd1)
) axi_crossbar (
	.clk(sys_clk),
	.m_axi_arready({cramsoc_dbus_ar_ready, cramsoc_axi_csr_ar_ready, cramsoc_dbus_peri_ar_ready}),
	.m_axi_awready({cramsoc_dbus_aw_ready, cramsoc_axi_csr_aw_ready, cramsoc_dbus_peri_aw_ready}),
	.m_axi_bid({cramsoc_dbus_b_param_id, cramsoc_axi_csr_b_param_id, cramsoc_dbus_peri_b_param_id}),
	.m_axi_bresp({cramsoc_dbus_b_payload_resp, cramsoc_axi_csr_b_payload_resp, cramsoc_dbus_peri_b_payload_resp}),
	.m_axi_buser({cramsoc_dbus_b_param_user, cramsoc_axi_csr_b_param_user, cramsoc_dbus_peri_b_param_user}),
	.m_axi_bvalid({cramsoc_dbus_b_valid, cramsoc_axi_csr_b_valid, cramsoc_dbus_peri_b_valid}),
	.m_axi_rdata({cramsoc_dbus_r_payload_data, cramsoc_axi_csr_r_payload_data, cramsoc_dbus_peri_r_payload_data}),
	.m_axi_rid({cramsoc_dbus_r_param_id, cramsoc_axi_csr_r_param_id, cramsoc_dbus_peri_r_param_id}),
	.m_axi_rlast({cramsoc_dbus_r_last, cramsoc_axi_csr_r_last, cramsoc_dbus_peri_r_last}),
	.m_axi_rresp({cramsoc_dbus_r_payload_resp, cramsoc_axi_csr_r_payload_resp, cramsoc_dbus_peri_r_payload_resp}),
	.m_axi_ruser({cramsoc_dbus_r_param_user, cramsoc_axi_csr_r_param_user, cramsoc_dbus_peri_r_param_user}),
	.m_axi_rvalid({cramsoc_dbus_r_valid, cramsoc_axi_csr_r_valid, cramsoc_dbus_peri_r_valid}),
	.m_axi_wready({cramsoc_dbus_w_ready, cramsoc_axi_csr_w_ready, cramsoc_dbus_peri_w_ready}),
	.rst(sys_rst),
	.s_axi_araddr({cramsoc_dbus_axi_ar_payload_addr}),
	.s_axi_arburst({cramsoc_dbus_axi_ar_payload_burst}),
	.s_axi_arcache({cramsoc_dbus_axi_ar_payload_cache}),
	.s_axi_arid({cramsoc_dbus_axi_ar_param_id}),
	.s_axi_arlen({cramsoc_dbus_axi_ar_payload_len}),
	.s_axi_arlock({cramsoc_dbus_axi_ar_payload_lock}),
	.s_axi_arprot({cramsoc_dbus_axi_ar_payload_prot}),
	.s_axi_arqos({cramsoc_dbus_axi_ar_payload_qos}),
	.s_axi_arsize({cramsoc_dbus_axi_ar_payload_size}),
	.s_axi_aruser({cramsoc_dbus_axi_ar_param_user}),
	.s_axi_arvalid({cramsoc_dbus_axi_ar_valid}),
	.s_axi_awaddr({cramsoc_dbus_axi_aw_payload_addr}),
	.s_axi_awburst({cramsoc_dbus_axi_aw_payload_burst}),
	.s_axi_awcache({cramsoc_dbus_axi_aw_payload_cache}),
	.s_axi_awid({cramsoc_dbus_axi_aw_param_id}),
	.s_axi_awlen({cramsoc_dbus_axi_aw_payload_len}),
	.s_axi_awlock({cramsoc_dbus_axi_aw_payload_lock}),
	.s_axi_awprot({cramsoc_dbus_axi_aw_payload_prot}),
	.s_axi_awqos({cramsoc_dbus_axi_aw_payload_qos}),
	.s_axi_awsize({cramsoc_dbus_axi_aw_payload_size}),
	.s_axi_awuser({cramsoc_dbus_axi_aw_param_user}),
	.s_axi_awvalid({cramsoc_dbus_axi_aw_valid}),
	.s_axi_bready({cramsoc_dbus_axi_b_ready}),
	.s_axi_rready({cramsoc_dbus_axi_r_ready}),
	.s_axi_wdata({cramsoc_dbus_axi_w_payload_data}),
	.s_axi_wlast({cramsoc_dbus_axi_w_last}),
	.s_axi_wstrb({cramsoc_dbus_axi_w_payload_strb}),
	.s_axi_wuser({cramsoc_dbus_axi_w_param_user}),
	.s_axi_wvalid({cramsoc_dbus_axi_w_valid}),
	.m_axi_araddr({cramsoc_dbus_ar_payload_addr, cramsoc_axi_csr_ar_payload_addr, cramsoc_dbus_peri_ar_payload_addr}),
	.m_axi_arburst({cramsoc_dbus_ar_payload_burst, cramsoc_axi_csr_ar_payload_burst, cramsoc_dbus_peri_ar_payload_burst}),
	.m_axi_arcache({cramsoc_dbus_ar_payload_cache, cramsoc_axi_csr_ar_payload_cache, cramsoc_dbus_peri_ar_payload_cache}),
	.m_axi_arid({cramsoc_dbus_ar_param_id, cramsoc_axi_csr_ar_param_id, cramsoc_dbus_peri_ar_param_id}),
	.m_axi_arlen({cramsoc_dbus_ar_payload_len, cramsoc_axi_csr_ar_payload_len, cramsoc_dbus_peri_ar_payload_len}),
	.m_axi_arlock({cramsoc_dbus_ar_payload_lock, cramsoc_axi_csr_ar_payload_lock, cramsoc_dbus_peri_ar_payload_lock}),
	.m_axi_arprot({cramsoc_dbus_ar_payload_prot, cramsoc_axi_csr_ar_payload_prot, cramsoc_dbus_peri_ar_payload_prot}),
	.m_axi_arqos({cramsoc_dbus_ar_payload_qos, cramsoc_axi_csr_ar_payload_qos, cramsoc_dbus_peri_ar_payload_qos}),
	.m_axi_arregion({cramsoc_dbus_ar_payload_region, cramsoc_axi_csr_ar_payload_region, cramsoc_dbus_peri_ar_payload_region}),
	.m_axi_arsize({cramsoc_dbus_ar_payload_size, cramsoc_axi_csr_ar_payload_size, cramsoc_dbus_peri_ar_payload_size}),
	.m_axi_aruser({cramsoc_dbus_ar_param_user, cramsoc_axi_csr_ar_param_user, cramsoc_dbus_peri_ar_param_user}),
	.m_axi_arvalid({cramsoc_dbus_ar_valid, cramsoc_axi_csr_ar_valid, cramsoc_dbus_peri_ar_valid}),
	.m_axi_awaddr({cramsoc_dbus_aw_payload_addr, cramsoc_axi_csr_aw_payload_addr, cramsoc_dbus_peri_aw_payload_addr}),
	.m_axi_awburst({cramsoc_dbus_aw_payload_burst, cramsoc_axi_csr_aw_payload_burst, cramsoc_dbus_peri_aw_payload_burst}),
	.m_axi_awcache({cramsoc_dbus_aw_payload_cache, cramsoc_axi_csr_aw_payload_cache, cramsoc_dbus_peri_aw_payload_cache}),
	.m_axi_awid({cramsoc_dbus_aw_param_id, cramsoc_axi_csr_aw_param_id, cramsoc_dbus_peri_aw_param_id}),
	.m_axi_awlen({cramsoc_dbus_aw_payload_len, cramsoc_axi_csr_aw_payload_len, cramsoc_dbus_peri_aw_payload_len}),
	.m_axi_awlock({cramsoc_dbus_aw_payload_lock, cramsoc_axi_csr_aw_payload_lock, cramsoc_dbus_peri_aw_payload_lock}),
	.m_axi_awprot({cramsoc_dbus_aw_payload_prot, cramsoc_axi_csr_aw_payload_prot, cramsoc_dbus_peri_aw_payload_prot}),
	.m_axi_awqos({cramsoc_dbus_aw_payload_qos, cramsoc_axi_csr_aw_payload_qos, cramsoc_dbus_peri_aw_payload_qos}),
	.m_axi_awregion({cramsoc_dbus_aw_payload_region, cramsoc_axi_csr_aw_payload_region, cramsoc_dbus_peri_aw_payload_region}),
	.m_axi_awsize({cramsoc_dbus_aw_payload_size, cramsoc_axi_csr_aw_payload_size, cramsoc_dbus_peri_aw_payload_size}),
	.m_axi_awuser({cramsoc_dbus_aw_param_user, cramsoc_axi_csr_aw_param_user, cramsoc_dbus_peri_aw_param_user}),
	.m_axi_awvalid({cramsoc_dbus_aw_valid, cramsoc_axi_csr_aw_valid, cramsoc_dbus_peri_aw_valid}),
	.m_axi_bready({cramsoc_dbus_b_ready, cramsoc_axi_csr_b_ready, cramsoc_dbus_peri_b_ready}),
	.m_axi_rready({cramsoc_dbus_r_ready, cramsoc_axi_csr_r_ready, cramsoc_dbus_peri_r_ready}),
	.m_axi_wdata({cramsoc_dbus_w_payload_data, cramsoc_axi_csr_w_payload_data, cramsoc_dbus_peri_w_payload_data}),
	.m_axi_wlast({cramsoc_dbus_w_last, cramsoc_axi_csr_w_last, cramsoc_dbus_peri_w_last}),
	.m_axi_wstrb({cramsoc_dbus_w_payload_strb, cramsoc_axi_csr_w_payload_strb, cramsoc_dbus_peri_w_payload_strb}),
	.m_axi_wuser({cramsoc_dbus_w_param_user, cramsoc_axi_csr_w_param_user, cramsoc_dbus_peri_w_param_user}),
	.m_axi_wvalid({cramsoc_dbus_w_valid, cramsoc_axi_csr_w_valid, cramsoc_dbus_peri_w_valid}),
	.s_axi_arready({cramsoc_dbus_axi_ar_ready}),
	.s_axi_awready({cramsoc_dbus_axi_aw_ready}),
	.s_axi_bid({cramsoc_dbus_axi_b_param_id}),
	.s_axi_bresp({cramsoc_dbus_axi_b_payload_resp}),
	.s_axi_buser({cramsoc_dbus_axi_b_param_user}),
	.s_axi_bvalid({cramsoc_dbus_axi_b_valid}),
	.s_axi_rdata({cramsoc_dbus_axi_r_payload_data}),
	.s_axi_rid({cramsoc_dbus_axi_r_param_id}),
	.s_axi_rlast({cramsoc_dbus_axi_r_last}),
	.s_axi_rresp({cramsoc_dbus_axi_r_payload_resp}),
	.s_axi_ruser({cramsoc_dbus_axi_r_param_user}),
	.s_axi_rvalid({cramsoc_dbus_axi_r_valid}),
	.s_axi_wready({cramsoc_dbus_axi_w_ready})
);

VexRiscvAxi4 VexRiscvAxi4(
		.rbif_rdram1kx32		(rbif_rdram1kx32[2:5]),
		.rbif_rdram128x22		(rbif_rdram128x22[0:7]),
		.rbif_rdram512x64		(rbif_rdram512x64[0:3]),
	.CMATPG(cramsoc_cmatpg),
	.CMBIST(cramsoc_cmbist),
	.clk(sys_clk),
	.dBusAxi_ar_ready(cramsoc_dbus_axi_ar_ready),
	.dBusAxi_aw_ready(cramsoc_dbus_axi_aw_ready),
	.dBusAxi_b_payload_id(cramsoc_dbus_axi_b_param_id),
	.dBusAxi_b_payload_resp(cramsoc_dbus_axi_b_payload_resp),
	.dBusAxi_b_valid(cramsoc_dbus_axi_b_valid),
	.dBusAxi_r_payload_data(cramsoc_dbus_axi_r_payload_data),
	.dBusAxi_r_payload_id(cramsoc_dbus_axi_r_param_id),
	.dBusAxi_r_payload_last(cramsoc_dbus_axi_r_last),
	.dBusAxi_r_payload_resp(cramsoc_dbus_axi_r_payload_resp),
	.dBusAxi_r_valid(cramsoc_dbus_axi_r_valid),
	.dBusAxi_w_ready(cramsoc_dbus_axi_w_ready),
	.debugReset((~jtag_trst_n)),
	.externalInterruptArray(cramsoc_interrupt),
	.externalResetVector(cramsoc_vexriscvaxi_reset_mux),
	.iBusAxi_ar_ready(cramsoc_ibus_axi_ar_ready),
	.iBusAxi_r_payload_data(cramsoc_ibus_axi_r_payload_data),
	.iBusAxi_r_payload_id(cramsoc_ibus_axi_r_param_id),
	.iBusAxi_r_payload_last(cramsoc_ibus_axi_r_last),
	.iBusAxi_r_payload_resp(cramsoc_ibus_axi_r_payload_resp),
	.iBusAxi_r_valid(cramsoc_ibus_axi_r_valid),
	.jtag_tck(jtag_tck),
	.jtag_tdi(jtag_tdi),
	.jtag_tms(jtag_tms),
	.reset((sys_rst | debug_reset)),
	.softwareInterrupt(1'd0),
	.sramtrm(cramsoc_vexsramtrm),
	.timerInterrupt(1'd0),
	.CsrPlugin_inWfi(cramsoc_wfi_active),
	.CsrPlugin_privilege(cramsoc_privilege),
	.MmuPlugin_satp_asid(cramsoc_satp_asid),
	.MmuPlugin_satp_mode(cramsoc_satp_mode),
	.MmuPlugin_satp_ppn(cramsoc_satp_ppn),
	.dBusAxi_ar_payload_addr(cramsoc_dbus_axi_ar_payload_addr),
	.dBusAxi_ar_payload_burst(cramsoc_dbus_axi_ar_payload_burst),
	.dBusAxi_ar_payload_cache(cramsoc_dbus_axi_ar_payload_cache),
	.dBusAxi_ar_payload_id(cramsoc_dbus_axi_ar_param_id),
	.dBusAxi_ar_payload_len(cramsoc_dbus_axi_ar_payload_len),
	.dBusAxi_ar_payload_lock(cramsoc_dbus_axi_ar_payload_lock),
	.dBusAxi_ar_payload_prot(cramsoc_dbus_axi_ar_payload_prot),
	.dBusAxi_ar_payload_qos(cramsoc_dbus_axi_ar_payload_qos),
	.dBusAxi_ar_payload_region(cramsoc_dbus_axi_ar_payload_region),
	.dBusAxi_ar_payload_size(cramsoc_dbus_axi_ar_payload_size),
	.dBusAxi_ar_valid(cramsoc_dbus_axi_ar_valid),
	.dBusAxi_aw_payload_addr(cramsoc_dbus_axi_aw_payload_addr),
	.dBusAxi_aw_payload_burst(cramsoc_dbus_axi_aw_payload_burst),
	.dBusAxi_aw_payload_cache(cramsoc_dbus_axi_aw_payload_cache),
	.dBusAxi_aw_payload_id(cramsoc_dbus_axi_aw_param_id),
	.dBusAxi_aw_payload_len(cramsoc_dbus_axi_aw_payload_len),
	.dBusAxi_aw_payload_lock(cramsoc_dbus_axi_aw_payload_lock),
	.dBusAxi_aw_payload_prot(cramsoc_dbus_axi_aw_payload_prot),
	.dBusAxi_aw_payload_qos(cramsoc_dbus_axi_aw_payload_qos),
	.dBusAxi_aw_payload_region(cramsoc_dbus_axi_aw_payload_region),
	.dBusAxi_aw_payload_size(cramsoc_dbus_axi_aw_payload_size),
	.dBusAxi_aw_valid(cramsoc_dbus_axi_aw_valid),
	.dBusAxi_b_ready(cramsoc_dbus_axi_b_ready),
	.dBusAxi_r_ready(cramsoc_dbus_axi_r_ready),
	.dBusAxi_w_payload_data(cramsoc_dbus_axi_w_payload_data),
	.dBusAxi_w_payload_last(cramsoc_dbus_axi_w_last),
	.dBusAxi_w_payload_strb(cramsoc_dbus_axi_w_payload_strb),
	.dBusAxi_w_valid(cramsoc_dbus_axi_w_valid),
	.debug_resetOut(o_resetOut),
	.iBusAxi_ar_payload_addr(cramsoc_ibus_axi_ar_payload_addr),
	.iBusAxi_ar_payload_burst(cramsoc_ibus_axi_ar_payload_burst),
	.iBusAxi_ar_payload_cache(cramsoc_ibus_axi_ar_payload_cache),
	.iBusAxi_ar_payload_id(cramsoc_ibus_axi_ar_param_id),
	.iBusAxi_ar_payload_len(cramsoc_ibus_axi_ar_payload_len),
	.iBusAxi_ar_payload_lock(cramsoc_ibus_axi_ar_payload_lock),
	.iBusAxi_ar_payload_prot(cramsoc_ibus_axi_ar_payload_prot),
	.iBusAxi_ar_payload_qos(cramsoc_ibus_axi_ar_payload_qos),
	.iBusAxi_ar_payload_region(cramsoc_ibus_axi_ar_payload_region),
	.iBusAxi_ar_payload_size(cramsoc_ibus_axi_ar_payload_size),
	.iBusAxi_ar_valid(cramsoc_ibus_axi_ar_valid),
	.iBusAxi_r_ready(cramsoc_ibus_axi_r_ready),
	.jtag_tdo(jtag_tdo)
);

endmodule

// -----------------------------------------------------------------------------
//  Auto-Generated by LiteX on 2025-02-08 04:21:33.
//------------------------------------------------------------------------------
