// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

// -----------------------------------------------------------------------------
// Auto-Generated by:        __   _ __      _  __
//                          / /  (_) /____ | |/_/
//                         / /__/ / __/ -_)>  <
//                        /____/_/\__/\__/_/|_|
//                     Build your hardware, easily!
//                   https://github.com/enjoy-digital/litex
//
// Filename   : bio_tb.v
// Device     : generic
// LiteX sha1 : 5375731c
// Date       : 2024-11-22 15:27:29
//------------------------------------------------------------------------------

`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// Module
//------------------------------------------------------------------------------

module bio_tb (
    input  wire          sim_trace,
    input  wire          reset,
    input  wire          clk,
    input  wire   [31:0] test,
    inout  wire   [31:0] gpio
);


//------------------------------------------------------------------------------
// Signals
//------------------------------------------------------------------------------

wire          sys_clk;
wire          sys_rst;
wire          i2c;
wire          force_1;
wire   [15:0] force_val;
reg           i2c_scl = 1'd0;
reg           i2c_sda = 1'd0;
reg           i2c_scl_d = 1'd0;
reg           i2c_sda_d = 1'd0;
reg     [3:0] i2c_ctr = 4'd0;
reg     [7:0] i2c_adr_in = 8'd0;
reg     [7:0] i2c_dout = 8'd0;
reg           zero = 1'd0;
reg           i2c_sda_controller_drive_low = 1'd0;
reg           i2c_sda_peripheral_drive_low = 1'd0;
reg    [31:0] gpio_o = 32'd0;
reg    [31:0] gpio_i = 32'd0;
reg    [31:0] gpio_oe = 32'd0;
wire          tstriple0_o;
wire          tstriple0_oe;
wire          tstriple0_i;
wire          tstriple1_o;
wire          tstriple1_oe;
wire          tstriple1_i;
wire          tstriple2_o;
wire          tstriple2_oe;
wire          tstriple2_i;
wire          tstriple3_o;
wire          tstriple3_oe;
wire          tstriple3_i;
wire          tstriple4_o;
wire          tstriple4_oe;
wire          tstriple4_i;
wire          tstriple5_o;
wire          tstriple5_oe;
wire          tstriple5_i;
wire          tstriple6_o;
wire          tstriple6_oe;
wire          tstriple6_i;
wire          tstriple7_o;
wire          tstriple7_oe;
wire          tstriple7_i;
wire          tstriple8_o;
wire          tstriple8_oe;
wire          tstriple8_i;
wire          tstriple9_o;
wire          tstriple9_oe;
wire          tstriple9_i;
wire          tstriple10_o;
wire          tstriple10_oe;
wire          tstriple10_i;
wire          tstriple11_o;
wire          tstriple11_oe;
wire          tstriple11_i;
wire          tstriple12_o;
wire          tstriple12_oe;
wire          tstriple12_i;
wire          tstriple13_o;
wire          tstriple13_oe;
wire          tstriple13_i;
wire          tstriple14_o;
wire          tstriple14_oe;
wire          tstriple14_i;
wire          tstriple15_o;
wire          tstriple15_oe;
wire          tstriple15_i;
wire          tstriple16_o;
wire          tstriple16_oe;
wire          tstriple16_i;
wire          tstriple17_o;
wire          tstriple17_oe;
wire          tstriple17_i;
wire          tstriple18_o;
wire          tstriple18_oe;
wire          tstriple18_i;
wire          tstriple19_o;
wire          tstriple19_oe;
wire          tstriple19_i;
wire          tstriple20_o;
wire          tstriple20_oe;
wire          tstriple20_i;
wire          tstriple21_o;
wire          tstriple21_oe;
wire          tstriple21_i;
wire          tstriple22_o;
wire          tstriple22_oe;
wire          tstriple22_i;
wire          tstriple23_o;
wire          tstriple23_oe;
wire          tstriple23_i;
wire          tstriple24_o;
wire          tstriple24_oe;
wire          tstriple24_i;
wire          tstriple25_o;
wire          tstriple25_oe;
wire          tstriple25_i;
wire          tstriple26_o;
wire          tstriple26_oe;
wire          tstriple26_i;
wire          tstriple27_o;
wire          tstriple27_oe;
wire          tstriple27_i;
wire          tstriple28_o;
wire          tstriple28_oe;
wire          tstriple28_i;
wire          tstriple29_o;
wire          tstriple29_oe;
wire          tstriple29_i;
wire          tstriple30_o;
wire          tstriple30_oe;
wire          tstriple30_i;
wire          tstriple31_o;
wire          tstriple31_oe;
wire          tstriple31_i;
reg     [2:0] state = 3'd0;
reg     [2:0] next_state = 3'd0;
reg     [3:0] i2c_ctr_next_value = 4'd0;
reg           i2c_ctr_next_value_ce = 1'd0;
reg     [7:0] i2c_adr_in_f_next_value = 8'd0;
reg           i2c_adr_in_f_next_value_ce = 1'd0;
reg     [7:0] i2c_dout_t_next_value = 8'd0;
reg           i2c_dout_t_next_value_ce = 1'd0;

//------------------------------------------------------------------------------
// Combinatorial Logic
//------------------------------------------------------------------------------

assign sys_clk = clk;
assign sys_rst = reset;
assign i2c = test[0];
assign force_1 = test[1];
assign force_val = test[31:16];
assign tstriple0_oe = gpio_oe[0];
assign tstriple0_o = gpio_o[0];
assign tstriple1_oe = gpio_oe[1];
assign tstriple1_o = gpio_o[1];
assign tstriple2_oe = gpio_oe[2];
assign tstriple2_o = gpio_o[2];
assign tstriple3_oe = gpio_oe[3];
assign tstriple3_o = gpio_o[3];
assign tstriple4_oe = gpio_oe[4];
assign tstriple4_o = gpio_o[4];
assign tstriple5_oe = gpio_oe[5];
assign tstriple5_o = gpio_o[5];
assign tstriple6_oe = gpio_oe[6];
assign tstriple6_o = gpio_o[6];
assign tstriple7_oe = gpio_oe[7];
assign tstriple7_o = gpio_o[7];
assign tstriple8_oe = gpio_oe[8];
assign tstriple8_o = gpio_o[8];
assign tstriple9_oe = gpio_oe[9];
assign tstriple9_o = gpio_o[9];
assign tstriple10_oe = gpio_oe[10];
assign tstriple10_o = gpio_o[10];
assign tstriple11_oe = gpio_oe[11];
assign tstriple11_o = gpio_o[11];
assign tstriple12_oe = gpio_oe[12];
assign tstriple12_o = gpio_o[12];
assign tstriple13_oe = gpio_oe[13];
assign tstriple13_o = gpio_o[13];
assign tstriple14_oe = gpio_oe[14];
assign tstriple14_o = gpio_o[14];
assign tstriple15_oe = gpio_oe[15];
assign tstriple15_o = gpio_o[15];
assign tstriple16_oe = gpio_oe[16];
assign tstriple16_o = gpio_o[16];
assign tstriple17_oe = gpio_oe[17];
assign tstriple17_o = gpio_o[17];
assign tstriple18_oe = gpio_oe[18];
assign tstriple18_o = gpio_o[18];
assign tstriple19_oe = gpio_oe[19];
assign tstriple19_o = gpio_o[19];
assign tstriple20_oe = gpio_oe[20];
assign tstriple20_o = gpio_o[20];
assign tstriple21_oe = gpio_oe[21];
assign tstriple21_o = gpio_o[21];
assign tstriple22_oe = gpio_oe[22];
assign tstriple22_o = gpio_o[22];
assign tstriple23_oe = gpio_oe[23];
assign tstriple23_o = gpio_o[23];
assign tstriple24_oe = gpio_oe[24];
assign tstriple24_o = gpio_o[24];
assign tstriple25_oe = gpio_oe[25];
assign tstriple25_o = gpio_o[25];
assign tstriple26_oe = gpio_oe[26];
assign tstriple26_o = gpio_o[26];
assign tstriple27_oe = gpio_oe[27];
assign tstriple27_o = gpio_o[27];
assign tstriple28_oe = gpio_oe[28];
assign tstriple28_o = gpio_o[28];
assign tstriple29_oe = gpio_oe[29];
assign tstriple29_o = gpio_o[29];
assign tstriple30_oe = gpio_oe[30];
assign tstriple30_o = gpio_o[30];
always @(*) begin
    gpio_i <= 32'd0;
    gpio_i[0] <= tstriple0_i;
    gpio_i[1] <= tstriple1_i;
    gpio_i[2] <= tstriple2_i;
    gpio_i[3] <= tstriple3_i;
    gpio_i[4] <= tstriple4_i;
    gpio_i[5] <= tstriple5_i;
    gpio_i[6] <= tstriple6_i;
    gpio_i[7] <= tstriple7_i;
    gpio_i[8] <= tstriple8_i;
    gpio_i[9] <= tstriple9_i;
    gpio_i[10] <= tstriple10_i;
    gpio_i[11] <= tstriple11_i;
    gpio_i[12] <= tstriple12_i;
    gpio_i[13] <= tstriple13_i;
    gpio_i[14] <= tstriple14_i;
    gpio_i[15] <= tstriple15_i;
    gpio_i[16] <= tstriple16_i;
    gpio_i[17] <= tstriple17_i;
    gpio_i[18] <= tstriple18_i;
    gpio_i[19] <= tstriple19_i;
    gpio_i[20] <= tstriple20_i;
    gpio_i[21] <= tstriple21_i;
    gpio_i[22] <= tstriple22_i;
    gpio_i[23] <= tstriple23_i;
    gpio_i[24] <= tstriple24_i;
    gpio_i[25] <= tstriple25_i;
    gpio_i[26] <= tstriple26_i;
    gpio_i[27] <= tstriple27_i;
    gpio_i[28] <= tstriple28_i;
    gpio_i[29] <= tstriple29_i;
    gpio_i[30] <= tstriple30_i;
    gpio_i[31] <= tstriple31_i;
end
assign tstriple31_oe = gpio_oe[31];
assign tstriple31_o = gpio_o[31];
always @(*) begin
    gpio_oe <= 32'd0;
    i2c_scl <= 1'd0;
    i2c_sda <= 1'd0;
    gpio_o <= 32'd0;
    if (force_1) begin
        gpio_o[0] <= force_val[0];
        gpio_oe[0] <= 1'd1;
    end else begin
        gpio_oe[0] <= 1'd0;
        gpio_o[0] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[1] <= force_val[1];
        gpio_oe[1] <= 1'd1;
    end else begin
        gpio_oe[1] <= 1'd0;
        gpio_o[1] <= 1'd0;
    end
    if (i2c) begin
        i2c_sda <= gpio_i[2];
        gpio_o[2] <= 1'd0;
        gpio_oe[2] <= (i2c_sda_controller_drive_low | i2c_sda_peripheral_drive_low);
    end else begin
        if (force_1) begin
            gpio_oe[2] <= 1'd1;
            gpio_o[2] <= force_val[2];
        end else begin
            gpio_oe[2] <= 1'd0;
        end
    end
    if (i2c) begin
        i2c_scl <= gpio_i[3];
    end else begin
        if (force_1) begin
            gpio_o[3] <= force_val[3];
            gpio_oe[3] <= 1'd1;
        end else begin
            gpio_oe[3] <= 1'd0;
        end
    end
    if (force_1) begin
        gpio_o[4] <= force_val[4];
        gpio_oe[4] <= 1'd1;
    end else begin
        gpio_oe[4] <= 1'd0;
        gpio_o[4] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[5] <= force_val[5];
        gpio_oe[5] <= 1'd1;
    end else begin
        gpio_oe[5] <= 1'd0;
        gpio_o[5] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[6] <= force_val[6];
        gpio_oe[6] <= 1'd1;
    end else begin
        gpio_oe[6] <= 1'd0;
        gpio_o[6] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[7] <= force_val[7];
        gpio_oe[7] <= 1'd1;
    end else begin
        gpio_oe[7] <= 1'd0;
        gpio_o[7] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[8] <= force_val[8];
        gpio_oe[8] <= 1'd1;
    end else begin
        gpio_oe[8] <= 1'd0;
        gpio_o[8] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[9] <= force_val[9];
        gpio_oe[9] <= 1'd1;
    end else begin
        gpio_oe[9] <= 1'd0;
        gpio_o[9] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[10] <= force_val[10];
        gpio_oe[10] <= 1'd1;
    end else begin
        gpio_oe[10] <= 1'd0;
        gpio_o[10] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[11] <= force_val[11];
        gpio_oe[11] <= 1'd1;
    end else begin
        gpio_oe[11] <= 1'd0;
        gpio_o[11] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[12] <= force_val[12];
        gpio_oe[12] <= 1'd1;
    end else begin
        gpio_oe[12] <= 1'd0;
        gpio_o[12] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[13] <= force_val[13];
        gpio_oe[13] <= 1'd1;
    end else begin
        gpio_oe[13] <= 1'd0;
        gpio_o[13] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[14] <= force_val[14];
        gpio_oe[14] <= 1'd1;
    end else begin
        gpio_oe[14] <= 1'd0;
        gpio_o[14] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[15] <= force_val[15];
        gpio_oe[15] <= 1'd1;
    end else begin
        gpio_oe[15] <= 1'd0;
        gpio_o[15] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[16] <= (~force_val[0]);
        gpio_oe[16] <= 1'd1;
    end else begin
        gpio_oe[16] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[17] <= (~force_val[1]);
        gpio_oe[17] <= 1'd1;
    end else begin
        gpio_oe[17] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[18] <= (~force_val[2]);
        gpio_oe[18] <= 1'd1;
    end else begin
        gpio_oe[18] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[19] <= (~force_val[3]);
        gpio_oe[19] <= 1'd1;
    end else begin
        gpio_oe[19] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[20] <= (~force_val[4]);
        gpio_oe[20] <= 1'd1;
    end else begin
        gpio_oe[20] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[21] <= (~force_val[5]);
        gpio_oe[21] <= 1'd1;
    end else begin
        gpio_oe[21] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[22] <= (~force_val[6]);
        gpio_oe[22] <= 1'd1;
    end else begin
        gpio_oe[22] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[23] <= (~force_val[7]);
        gpio_oe[23] <= 1'd1;
    end else begin
        gpio_oe[23] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[24] <= (~force_val[8]);
        gpio_oe[24] <= 1'd1;
    end else begin
        gpio_oe[24] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[25] <= (~force_val[9]);
        gpio_oe[25] <= 1'd1;
    end else begin
        gpio_oe[25] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[26] <= (~force_val[10]);
        gpio_oe[26] <= 1'd1;
    end else begin
        gpio_oe[26] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[27] <= (~force_val[11]);
        gpio_oe[27] <= 1'd1;
    end else begin
        gpio_oe[27] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[28] <= (~force_val[12]);
        gpio_oe[28] <= 1'd1;
    end else begin
        gpio_oe[28] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[29] <= (~force_val[13]);
        gpio_oe[29] <= 1'd1;
    end else begin
        gpio_oe[29] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[30] <= (~force_val[14]);
        gpio_oe[30] <= 1'd1;
    end else begin
        gpio_oe[30] <= 1'd0;
    end
    if (force_1) begin
        gpio_o[31] <= (~force_val[15]);
        gpio_oe[31] <= 1'd1;
    end else begin
        gpio_oe[31] <= 1'd0;
    end
end
always @(*) begin
    i2c_adr_in_f_next_value <= 8'd0;
    i2c_adr_in_f_next_value_ce <= 1'd0;
    next_state <= 3'd0;
    i2c_sda_controller_drive_low <= 1'd0;
    i2c_sda_peripheral_drive_low <= 1'd0;
    i2c_ctr_next_value <= 4'd0;
    i2c_ctr_next_value_ce <= 1'd0;
    i2c_dout_t_next_value <= 8'd0;
    i2c_dout_t_next_value_ce <= 1'd0;
    next_state <= state;
    case (state)
        1'd1: begin
            if ((((i2c_sda_d & (~i2c_sda)) & i2c_scl) & i2c_scl_d)) begin
                i2c_ctr_next_value <= 4'd8;
                i2c_ctr_next_value_ce <= 1'd1;
                next_state <= 1'd1;
            end else begin
                if (((((~i2c_sda_d) & i2c_sda) & i2c_scl) & i2c_scl_d)) begin
                    next_state <= 1'd0;
                end else begin
                    if ((i2c_scl & (~i2c_scl_d))) begin
                        i2c_ctr_next_value <= (i2c_ctr - 1'd1);
                        i2c_ctr_next_value_ce <= 1'd1;
                        if ((i2c_ctr != 1'd0)) begin
                            i2c_adr_in_f_next_value <= {i2c_adr_in[6:0], i2c_sda};
                            i2c_adr_in_f_next_value_ce <= 1'd1;
                        end
                    end else begin
                        if (((~i2c_scl) & i2c_scl_d)) begin
                            if ((i2c_ctr == 1'd0)) begin
                                next_state <= 2'd2;
                            end
                        end
                    end
                end
            end
        end
        2'd2: begin
            if ((i2c_adr_in != 5'd23)) begin
                i2c_sda_peripheral_drive_low <= 1'd1;
            end
            if (((((~i2c_sda_d) & i2c_sda) & i2c_scl) & i2c_scl_d)) begin
                next_state <= 1'd0;
            end else begin
                if (((~i2c_scl) & i2c_scl_d)) begin
                    i2c_dout_t_next_value <= (~i2c_adr_in);
                    i2c_dout_t_next_value_ce <= 1'd1;
                    if ((i2c_adr_in != 5'd23)) begin
                        i2c_ctr_next_value <= 4'd8;
                        i2c_ctr_next_value_ce <= 1'd1;
                        if (i2c_adr_in[0]) begin
                            next_state <= 2'd3;
                        end else begin
                            next_state <= 1'd1;
                        end
                    end else begin
                        next_state <= 1'd0;
                    end
                end
            end
        end
        2'd3: begin
            if (((((~i2c_sda_d) & i2c_sda) & i2c_scl) & i2c_scl_d)) begin
                next_state <= 1'd0;
            end else begin
                if (((~i2c_scl) & i2c_scl_d)) begin
                    i2c_ctr_next_value <= (i2c_ctr - 1'd1);
                    i2c_ctr_next_value_ce <= 1'd1;
                    if ((i2c_ctr != 1'd0)) begin
                        i2c_dout_t_next_value <= {i2c_dout[6:0], zero};
                        i2c_dout_t_next_value_ce <= 1'd1;
                    end
                end else begin
                    if ((i2c_scl & (~i2c_scl_d))) begin
                        if ((i2c_ctr == 1'd0)) begin
                            next_state <= 3'd4;
                        end
                    end
                end
            end
            i2c_sda_controller_drive_low <= (~i2c_dout[7]);
        end
        3'd4: begin
            if (((((~i2c_sda_d) & i2c_sda) & i2c_scl) & i2c_scl_d)) begin
                next_state <= 1'd0;
            end else begin
                if (((~i2c_scl) & i2c_scl_d)) begin
                    next_state <= 1'd0;
                end
            end
        end
        default: begin
            if ((((i2c_sda_d & (~i2c_sda)) & i2c_scl) & i2c_scl_d)) begin
                i2c_ctr_next_value <= 4'd8;
                i2c_ctr_next_value_ce <= 1'd1;
                next_state <= 1'd1;
            end
        end
    endcase
end


//------------------------------------------------------------------------------
// Synchronous Logic
//------------------------------------------------------------------------------

always @(posedge sys_clk) begin
    i2c_sda_d <= i2c_sda;
    i2c_scl_d <= i2c_scl;
    state <= next_state;
    if (i2c_ctr_next_value_ce) begin
        i2c_ctr <= i2c_ctr_next_value;
    end
    if (i2c_adr_in_f_next_value_ce) begin
        i2c_adr_in <= i2c_adr_in_f_next_value;
    end
    if (i2c_dout_t_next_value_ce) begin
        i2c_dout <= i2c_dout_t_next_value;
    end
    if (sys_rst) begin
        i2c_scl_d <= 1'd0;
        i2c_sda_d <= 1'd0;
        i2c_ctr <= 4'd0;
        i2c_adr_in <= 8'd0;
        i2c_dout <= 8'd0;
        state <= 3'd0;
    end
end


//------------------------------------------------------------------------------
// Specialized Logic
//------------------------------------------------------------------------------

assign gpio[0] = tstriple0_oe ? tstriple0_o : 1'bz;
assign tstriple0_i = gpio[0];

assign gpio[1] = tstriple1_oe ? tstriple1_o : 1'bz;
assign tstriple1_i = gpio[1];

assign gpio[2] = tstriple2_oe ? tstriple2_o : 1'bz;
assign tstriple2_i = gpio[2];

assign gpio[3] = tstriple3_oe ? tstriple3_o : 1'bz;
assign tstriple3_i = gpio[3];

assign gpio[4] = tstriple4_oe ? tstriple4_o : 1'bz;
assign tstriple4_i = gpio[4];

assign gpio[5] = tstriple5_oe ? tstriple5_o : 1'bz;
assign tstriple5_i = gpio[5];

assign gpio[6] = tstriple6_oe ? tstriple6_o : 1'bz;
assign tstriple6_i = gpio[6];

assign gpio[7] = tstriple7_oe ? tstriple7_o : 1'bz;
assign tstriple7_i = gpio[7];

assign gpio[8] = tstriple8_oe ? tstriple8_o : 1'bz;
assign tstriple8_i = gpio[8];

assign gpio[9] = tstriple9_oe ? tstriple9_o : 1'bz;
assign tstriple9_i = gpio[9];

assign gpio[10] = tstriple10_oe ? tstriple10_o : 1'bz;
assign tstriple10_i = gpio[10];

assign gpio[11] = tstriple11_oe ? tstriple11_o : 1'bz;
assign tstriple11_i = gpio[11];

assign gpio[12] = tstriple12_oe ? tstriple12_o : 1'bz;
assign tstriple12_i = gpio[12];

assign gpio[13] = tstriple13_oe ? tstriple13_o : 1'bz;
assign tstriple13_i = gpio[13];

assign gpio[14] = tstriple14_oe ? tstriple14_o : 1'bz;
assign tstriple14_i = gpio[14];

assign gpio[15] = tstriple15_oe ? tstriple15_o : 1'bz;
assign tstriple15_i = gpio[15];

assign gpio[16] = tstriple16_oe ? tstriple16_o : 1'bz;
assign tstriple16_i = gpio[16];

assign gpio[17] = tstriple17_oe ? tstriple17_o : 1'bz;
assign tstriple17_i = gpio[17];

assign gpio[18] = tstriple18_oe ? tstriple18_o : 1'bz;
assign tstriple18_i = gpio[18];

assign gpio[19] = tstriple19_oe ? tstriple19_o : 1'bz;
assign tstriple19_i = gpio[19];

assign gpio[20] = tstriple20_oe ? tstriple20_o : 1'bz;
assign tstriple20_i = gpio[20];

assign gpio[21] = tstriple21_oe ? tstriple21_o : 1'bz;
assign tstriple21_i = gpio[21];

assign gpio[22] = tstriple22_oe ? tstriple22_o : 1'bz;
assign tstriple22_i = gpio[22];

assign gpio[23] = tstriple23_oe ? tstriple23_o : 1'bz;
assign tstriple23_i = gpio[23];

assign gpio[24] = tstriple24_oe ? tstriple24_o : 1'bz;
assign tstriple24_i = gpio[24];

assign gpio[25] = tstriple25_oe ? tstriple25_o : 1'bz;
assign tstriple25_i = gpio[25];

assign gpio[26] = tstriple26_oe ? tstriple26_o : 1'bz;
assign tstriple26_i = gpio[26];

assign gpio[27] = tstriple27_oe ? tstriple27_o : 1'bz;
assign tstriple27_i = gpio[27];

assign gpio[28] = tstriple28_oe ? tstriple28_o : 1'bz;
assign tstriple28_i = gpio[28];

assign gpio[29] = tstriple29_oe ? tstriple29_o : 1'bz;
assign tstriple29_i = gpio[29];

assign gpio[30] = tstriple30_oe ? tstriple30_o : 1'bz;
assign tstriple30_i = gpio[30];

assign gpio[31] = tstriple31_oe ? tstriple31_o : 1'bz;
assign tstriple31_i = gpio[31];

endmodule

// -----------------------------------------------------------------------------
//  Auto-Generated by LiteX on 2024-11-22 15:27:29.
//------------------------------------------------------------------------------
