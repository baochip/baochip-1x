// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/RtcApbif.v"
`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/RtcControl.v"
`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/RtcCounter.v"
`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/RtcInterrupt.v"
//`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/RtcParams.v"
`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/RtcRevAnd.v"
`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/RtcSynctoPCLK.v"
`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/RtcUpdate.v"
`include "ips/PL031_RTC/PL031-BU-01000-r1p3-00rel0/rtc_pl031/verilog/rtl_source/Rtc.v"
