// (c) Copyright 2024 CrossBar, Inc.
//
// SPDX-FileCopyrightText: 2024 CrossBar, Inc.
// SPDX-License-Identifier: CERN-OHL-W-2.0
//
// This documentation and source code is licensed under the CERN Open Hardware
// License Version 2 – Weakly Reciprocal (http://ohwr.org/cernohl; the
// “License”). Your use of any source code herein is governed by the License.
//
// You may redistribute and modify this documentation under the terms of the
// License. This documentation and source code is distributed WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTY, MERCHANTABILITY, SATISFACTORY QUALITY OR FITNESS FOR A
// PARTICULAR PURPOSE. Please see the License for the specific language governing
// permissions and limitations under the License.

`include "include/common_cell_inc.sv"

`include "modules/core/rtl/tcmram.sv"
`include "modules/core/rtl/cm7sys_tcm.sv"
`include "modules/core/rtl/cm7sys.sv"

`include "modules/core/rtl/itcm16kx18x2.sv"

`ifdef SIM
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_tcm_ram.v"

`define ARM_UD_MODEL
`define ARM_DISABLE_EMA_CHECK
`include "asic_top/lib/arm_sram_macro/ram32kx72/ram32kx72.v"
`include "asic_top/lib/arm_sram_macro/ram8kx72/ram8kx72.v"
`include "asic_top/lib/arm_sram_macro/rf1kx72_srm/rf1kx72.v"
`include "asic_top/lib/arm_sram_macro/rf256x27_srm/rf256x27.v"
`include "asic_top/lib/arm_sram_macro/rf512x39_srm/rf512x39.v"
`include "asic_top/lib/arm_sram_macro/rf128x31_srm/rf128x31.v"

`ifdef TCMSVT
//`include "lib/arm_sram_macro/dtcm8kx36/dtcm8kx36.v"
//`include "lib/arm_sram_macro/itcm32kx18/itcm32kx18.v"
`else
`include "asic_top/lib/arm_sram_macro/dtcm8kx36_srm/dtcm8kx36.v"
//`include "asic_top/lib/arm_sram_macro/itcm32kx18_srm/itcm32kx18.v"
`include "asic_top/lib/arm_sram_macro/itcm16kx18/itcm16kx18.v"

`endif
//`include "rtl/model/bit_ram.v"
`endif

`include "modules/model/rtl/cm7cell_clkgate.v"
`include "modules/model/rtl/cm7top_cache_rams_daric.v"

`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_atb_sync.v"
//`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_decl.v"
`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_trace_out.v"
`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu.v"
`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_formatter.v"
`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_trace_fifo.v"
`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_apb_if.v"
`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_trace_clk.v"
`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_atb_fifo.v"
`include "ips/cortexm7/logical/cm7tpiu/verilog/cm7tpiu_trace_sync.v"
`include "ips/cortexm7/logical/cm7stb/verilog/cm7stb_slot.v"
`include "ips/cortexm7/logical/cm7stb/verilog/cm7stb.v"
//`include "ips/cortexm7/logical/cm7stb/verilog/cm7stb_defs.v"
//`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_params.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu.v"
//`include "ips/cortexm7/logical/cm7core/verilog/cm7core_decl.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_swizzle_store.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7pfu.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_rf.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_sbitx.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_full_t32_pre.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_swizzle_load.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_au.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_div.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_clz.v"
//`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_ualdis.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_rbit.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_fpu_small_t32_post.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_fpu_full_t32_post.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_extract.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_predec.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_front_end.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_sat_dbl.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dp1_alu.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_shift.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_gen_sat.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_masksel.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dp0.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_undef_small.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_full_t16_pre.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_prog_flow.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_small_t16_post.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_iq.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7pfu_fifo.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_small_t32_post.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_full_t16_post.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_maskgen.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_etm_intf.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_full_t32_post.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_agu.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_lu.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7pfu_btac.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_mac.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_alu_simd_sat.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7core.v"
`include "ips/cortexm7/logical/cm7core/verilog/cm7dpu_dec_undef_full.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_miu.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_sq_half.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_tcm.v"
//`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_decl.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_sq.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_lsu.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_pfu.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_ahbs.v"
`include "ips/cortexm7/logical/cm7tcu/verilog/cm7tcu_sq_fifo.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_pend_cell.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_int_state.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_pend_tree_stage.v"
//`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_param.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_actv_tree.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_pend_tree.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_preempt.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_reg.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_actv_cell.v"
//`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_decl.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_ppb_intf.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_actv_tree_stage.v"
//`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_param_instan.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic.v"
`include "ips/cortexm7/logical/cm7nvic/verilog/cm7nvic_main.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7cell_cdc_and.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_pmu_sync_reset.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_rst_send_set.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7cell_dcreg.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_sw_cdc_capt_reset.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7cell_dcctl.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7cell_semi_sync_flop.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_pmu_sync_set.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7cell_sync.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_cdc_send_data.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_cdc_random.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7cell_dccm.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_cdc_and.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_cdc_send.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_cdc_send_addr.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_cdc_send_reset.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_sw_cdc_capt_sync.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_cdc_capt_sync.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_cdc_mux.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_pmu_cdc_send_reset.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_dap_cdc_capt_sync.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_rst_sync.v"
`include "ips/cortexm7/logical/models/cells/generic/cm7_cdc_connect.v"
`include "ips/cortexm7/logical/cm7icu/verilog/cm7icu.v"
//`include "ips/cortexm7/logical/cm7icu/verilog/cm7icu_decl.v"
`include "ips/cortexm7/logical/cm7icu/verilog/cm7icu_ecc_check.v"
`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti_apb_if.v"
`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti_reg_p.v"
`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti_reg_c.v"
`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti_mapper.v"
`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti.v"
//`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti_constants.v"
`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti_ci.v"
//`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti_undefs.v"
`include "ips/cortexm7/logical/cm7cti/verilog/cm7cti_ti.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_sram.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_tcm_ram.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/CM7IKMCU.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_clk_gen.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_sys.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_misc_delay.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_ahb_interconnect.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_ahb_sram_bridge_64.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_rst_ctl.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_stclken_gen.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_ahb_rom_bridge.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_misc.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_ahb_gpio.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_rom.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_pmu.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/example_sys/cm7_ik_ahb_def_slv.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/cm7_ik_trace_capture.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/cm7_ik_poreset.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/cm7_ik_debug_driver.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/cm7_ik_clk_src.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/CORTEXM7INTEGRATIONCS_input_delay.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/cm7_ik_defs.v"
//`include "ips/cortexm7/logical/testbench/execution_tb/verilog/tbench.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7/tbench/cm7top_sys_cache_ram_test.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7/tbench/generic_functions.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7/tbench/generic_testprocess.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7/tbench/dummy_cm7top_clk.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7/tbench/CORTEXM7_cache_ram_testbench.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7TCM/tbench/example/generic/CM7_TCM_RAM.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7TCM/tbench/example/TCMLevel.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7TCM/tbench/generic_functions.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7TCM/tbench/generic_testprocess.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7TCM/tbench/CORTEXM7_tcm_ram_testbench.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7TCM/tbench/dummy_cm7top_clk.v"
//`include "ips/cortexm7/logical/testbench/ram_integration_tb/CORTEXM7TCM/tbench/cm7top_sys_tcm_ram_test.v"
`include "ips/cortexm7/logical/cm7lsu/verilog/cm7lsu.v"
//`include "ips/cortexm7/logical/cm7lsu/verilog/cm7lsu_decl.v"
`include "ips/cortexm7/logical/cm7lsu/verilog/cm7lsu_lsu.v"
`include "ips/cortexm7/logical/cm7lsu/verilog/cm7lsu_ahbp.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_hazarding.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_waddr_buf.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_linefill.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_axi_interface.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_write_arbiter.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_linefill_buffer.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_read_arbiter.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu.v"
//`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_decl.v"
`include "ips/cortexm7/logical/cm7biu/verilog/cm7biu_linefill_buffer_ev_fsm.v"
`include "ips/cortexm7/logical/cm7fpb/verilog/cm7fpb.v"
`include "ips/cortexm7/logical/cm7dcu/verilog/cm7dcu_utag_way.v"
`include "ips/cortexm7/logical/cm7dcu/verilog/cm7dcu_ecc_maint.v"
`include "ips/cortexm7/logical/cm7dcu/verilog/cm7dcu_cachearb.v"
//`include "ips/cortexm7/logical/cm7dcu/verilog/cm7dcu_defs.v"
`include "ips/cortexm7/logical/cm7dcu/verilog/cm7dcu.v"
`include "ips/cortexm7/logical/cm7dcu/verilog/cm7dcu_utag.v"
`include "ips/cortexm7/logical/cm7miu/verilog/cm7miu.v"
`include "ips/cortexm7/logical/cm7dwt/verilog/cm7dwt_if.v"
`include "ips/cortexm7/logical/cm7dwt/verilog/cm7dwt_comp_data.v"
`include "ips/cortexm7/logical/cm7dwt/verilog/cm7dwt.v"
`include "ips/cortexm7/logical/cm7dwt/verilog/cm7dwt_packet_gen_fifo.v"
`include "ips/cortexm7/logical/cm7dwt/verilog/cm7dwt_packet_gen.v"
`include "ips/cortexm7/logical/cm7dwt/verilog/cm7dwt_comp.v"
`include "ips/cortexm7/logical/cm7itm/verilog/cm7itm_arb.v"
`include "ips/cortexm7/logical/cm7itm/verilog/cm7itm_if.v"
`include "ips/cortexm7/logical/cm7itm/verilog/cm7itm_fifo_byte.v"
`include "ips/cortexm7/logical/cm7itm/verilog/cm7itm.v"
`include "ips/cortexm7/logical/cm7itm/verilog/cm7itm_emit.v"
`include "ips/cortexm7/logical/cm7itm/verilog/cm7itm_fifo.v"
`include "ips/cortexm7/logical/cm7itm/verilog/cm7itm_lts.v"
//`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_ap_mast_defs.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_dp.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_ap_mast.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_dp_jtag.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_dp_cdc.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_dp_pwr.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_ap.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_dp_sw.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_ap_cdc.v"
//`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_dp_sw_defs.v"
//`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_dp_jtag_defs.v"
`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_top.v"
//`include "ips/cortexm7/logical/cm7dap/verilog/cm7_dap_invariants.v"
`include "ips/cortexm7/logical/cm7dap/verilog/CM7DAP.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_generate32.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ext_ahbs.v"
////`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_decl_tcm_types.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dpu_dwt.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_repair32.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_pfu_icu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_eppb_ext.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_miu_tcu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_pfu_tcu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_lsu_ahbp.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_top_ext.v"
////`include "ips/cortexm7/logical/cortexm7/verilog/cm7_csetmm7_pc.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ext_miu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_check32.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_etm_ipipe.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_mpu_pfu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7aab_ahb_ext.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7top_clk.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ppb_slv.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_itm_ext.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dpu_trc.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/CORTEXM7.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_miu_dcu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_miu_icu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ppb_dcu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_tcu_tcm.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_fatal64.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_lsu_biu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_lsu_tcu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ppb_icu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7top_sys.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_icu_biu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_etm_dpipe.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dpu_icu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dwt_itm.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_lsu_stb.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_sva_liveness.v"
////`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_decl.v"
////`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_decl_types.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_pfu_ext.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dcu_biu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_icu_ram.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_axi_ext.v"
////`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_decl_ahb_types.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_stb_dpu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_lsu_stb_biu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_axi_tracker_writes.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ahbp_ext.v"
////`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ext_dc.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_repair64.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_nvic_dpu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_miu_biu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_fatal32.v"
////`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_defs.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dbg_atb.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ppb_tcu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_biu_ext.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_lsu_dcu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ahbd_dpu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dpu_ppb.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_generate64.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_ext_ahbd.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dpu_fpu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_stb_biu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dpu_pfu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dpu_lsu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_decl_axi_types.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_mpu_dpu.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dcu_stb.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_dcu_ram.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_check64.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_axi_tracker_reads.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_nvic_tcu.v"
`include "ips/cortexm7/logical/cm7ppb/verilog/cm7ppb.v"
`include "ips/cortexm7/logical/cm7ppb/verilog/cm7ppb_reg.v"
`include "ips/cortexm7/logical/cm7mpu/verilog/cm7mpu.v"

`include "ips/cortexm7/logical/cortexm7/verilog/cm7top_clk.v"
`include "ips/cortexm7/logical/cortexm7/verilog/cm7top_sys.v"

`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_generate32.v"
`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_repair32.v"
`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_check32.v"
`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_fatal64.v"
`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_repair64.v"
`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_fatal32.v"
`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_generate64.v"
`include "ips/cortexm7/logical/cortexm7/verilog/cortexm7_ecc_check64.v"
//`include "ips/cortexm7/logical/cortexm7/verilog/cm7_csetmm7_pc.v"


`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_div_quot_sel.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_cvt.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_div.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_gen_int_rounding.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_ctz_32.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_div.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_cvt.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_fpscr.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_clz_64.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_clz_24.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_alu.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_mask_gen.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_mask_gen.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_pack.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_unpack.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_reg_pipe.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_hp_unpack.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_alu.v"
//`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_params.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_round.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_mul.v"
//`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_decl.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_mul.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_hp_unpack.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_ctz_24.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_unpack.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_sp_add.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_round.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_shifter.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_gen_rounding.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_pack.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_clz_32.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_clz_pred_mult.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_rf.v"
`include "ips/cortexm7/logical/cm7fpu/verilog/cm7fpu_dp_add.v"

`include "ips/cortexm7/logical/models/cells/generic/DS02_multp_24.v"
`include "ips/cortexm7/logical/models/cells/generic/DS02_multp_32.v"


`include "ips/cortexm7/logical/cortexm7_integration/verilog/cm7_cs_apb_rom_table.v"
`include "ips/cortexm7/logical/cortexm7_integration/verilog/cm7_cs_apb_interconnect.v"
`include "ips/cortexm7/logical/cortexm7_integration/verilog/cm7_wic.v"
`include "ips/cortexm7/logical/cortexm7_integration/verilog/cm7_mcu_apb_interconnect.v"

//`include "ips/cortexm7/logical/cortexm7_integration/verilog/CORTEXM7INTEGRATIONCS_CONFIG.v"
`include "modules/core/rtl/CORTEXM7.v"
`include "modules/core/rtl/CORTEXM7INTEGRATIONCS.v"
//`include "ips/cortexm7/logical/cortexm7_integration/verilog/CORTEXM7INTEGRATIONMCU.v"
